�D�  d0 0 ��^ @_�_�-@ �       ��� ? ����
  @ 
      \�^ �_�_�� �       H� ����� @       h�^ ��_�� �       ��=  ��?�   �        ��^��_�� �       0�? ���?�	� � 	      ��^�a�_�` �       0�? ���?�	� �       ��^�!�_��0 �       ��? ��?�p �       ��^��_�   �       �?  ��?�� �       ��^��_�   �       � ���� @       ��~�@�� ` �        ��� =����
 @ 
      8�~ 7���� �       ��� + ���� @       �t~ ?,_��, �       |�� �?��� � @        |t~ �_�� � �        0�� ^ȿ���!� @ e      ��~ ?�� �       �� 4`���` @ +      p�^�/��_�� � 1      @� ����� @       ��^�A�_�P �       ��? @��?�@ �       p�^���_��� �       ��?  ��?�  �       P�^���_�� �       ��? ��?� �       p�^���_��� �       ��? 
 ��?�  �       `�^�	��_�� �       P�? 
���?�� �       x�^���_��� �       X�? ���?�� �       �^���_�� � 	      8�� 	������ @       X�~��_��� �       ��� @?��� x @       xt~ �_��� �       h�� �?���� @       �tz _�� �       � �� 8?���08 @ 8      �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            