���  d0 0 Hz, <�_�/�� �       � � ?P/�� P �        xz/�:��/�� �       � ��@���X �       � z/�@_�/�
� �       � �� /��   �        �z�Q_���� �       ` �� ����`� �        0z� �_���� �        � �� ������ �        �z� �_���� �        0 �� ����� �        �z�  _���8 �          �� ������ �        �z�  _���8 �        � ��U/���� �        �~
�� _�
��  �        � �}UP/��P �       � ~�����8 �@       � �
_��/�
_�� ��       � ~��W���� �T       � �UU �UU  ���      � ~ *� � *� ��U      z �   �/�   � ���      � ~ *��� *�� ��U      , �UU�/�UU� ���      �z������ �AP      X ���o��� ��       �z
���
�� �        � ��U�/���� �        �z��_��� �        � ��U ����� �        0z��_���� �        � ��@@����@ �        �z� q_���p �        P �� ������ �        �z� �_���� �        P �� ����U� �        hz� �_���� �        x �P �/��@� �        xz/� ��/��� �        � �@ h_�� x �        �~/� @?�/��� �        � �  �� �       �z.�@?�/�p �       � � @_��` �       (z> �?�?�!� � !      � � #_�� �       �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            