���  d0 0 ��> FCh�߹�Ch�߹�      ������ !
E���
      _���;ޠ
�'�0���?      M���e��,�%��,�%�:      k�����Ԁ B��[�C      �w����4� �u��      ��^��� �N��3?      7�S�y���%����-��      �?=?�l`���p�a�����      ;s�}����G笘�g[      ջ_?g*D����:t�ȱ�      ���?�� 8�?s%���      �|����� X �X<      ��_���I� ?�i� �      ����>?	��$ɚE��      ��x���'�T�'�TS      �����C 	�k�mP��      ����}(  S�l S�      :  ��Ŕ  )�׶  ��      �  �T�0\  9      Ҹ
�/@���/�  �      ~�W�������@ǀ  @      } �������   �      ; �������a�    �      ��~����A � [      ��� 4h?���Kl @ k      x�^�o��_�� �       X� :���� @       ��^�'A�_�@ �       ��? @��?�'@ � '      p�^���_� � �       ��?  ��?�  �       P�^���_�� �       ��?  ��?�  �       p�^���_�� �       ��?  ��?�  �       p�^���_�� �       P�? ���?�� �       x�^���_�� �       X�? ���?�� �       �^���_�� � 	      8�� 	������ @       X�~��_��� �       ��� @?��� h @       xt~ �_��� �       x�� �?���� @       �tz _�� �       � �� 8?���08 @ 8      �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            