�;� ld0 0 �!HP	@t!         �!HP	�x���(5wby      �}����k�Ɓ��      ��{�Η�|���F:Ԥ K      _���������L/� <Q:�      ����~�)  $�kH���P      i���� ɚ ݭ8� �"b      8ͺ���:�H �=a      �˴�?{�R����n���      �����΀1���xe�      �����"6=4Q�YƆ��       {����[DM�i3 �[��D      [�_��w���F*D�P      ��+��W��h7p9��Z      ���u?(��s#GP�=�X      o���Z�E��%a�x@8      �}��=c
d��@���      S����q7����*      �����# �bH      -��'MC�r4��0(*      G�r<��1�8���Vg0�      3�~����y�ۀ�V���>A      ������1@z�@&�g
       qf�w�e$�p2F G>f	(      eg�v;n"@kQ]I��P��      k��{���0N��      ^�ߘ�5�	���0���$      ������[#��<g3	      ��g3٫�a��T�=}�      ���}��&#���A�052      W>������%��]�j��x      ��{���i�5dc�1Ba      m��5Zo��0R0�9G      V��=2_&�QG0c?�     (�sO?�0�f
/!8�      #n9��&G��0 �      �&w �0�2D3d��0L~�   o  �2t �8au(�x�
?�   
  y� �����@�k�   v �� ���X_�	@���  �  ��X ��8���)x�? ti  L  x�� ^<_����ìGj ��� �  �� �U��.,�DP�m�  �  ^]� =^�'¡<�v�  >�  ?  =���o�M�&�Wm� >�  �� �x\���+��[?�� [  �� ������Bfo^@ E�  ݀ ������)$�7m` _�  ŀ ����ÃU�  ���׺��       wU�_�.����P� m�n��� �      =^���¡6X� v�?>~��       =�?�]o��M�&� Wm�����       ]xs�������s[ ?����[ �      }����݀��f o^M�E� �      �������)+� 7mo�_�        ������       7�sN���           