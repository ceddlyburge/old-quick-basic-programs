�;��fd0 0 �����  �� ��  �  ŀ ����k� ؉�X<� ;  ̀ ����#��=��s�  �  ?�� ���{P e�؄P�  �  e�� ��&a��b0EP�b0  0�  gq� o�&���4U��4  �  w�� o�2鏾� ��@A�(   � ��� _� ����|� �x   K ��� }�dXO��ihǠ  h m^L o�����L�� ��     �� &.��zY܄K���   �@�O�\�������     P����˾N*p� s-�C�     ��o�s��=z5�}��XE�      ���}�� ��s�O�}`�      o�������Ʒa��aC8      ���ǿc}:d��@�#�X      S�;����|w����*      ������>�� !bH      -�?��MC�s4��0(*      G�s<��1�9���Vg0�      3�����y�ۀ�V���>A      ������1@z�@&�g       qf�w�e%�p2F E<f(      ee�v3n#�kY]H�P��      k��{����0N�C��      ^�_��5�)���0���$      ������!~��g3	      ��g3٨J
a��Tc=m�      �Zk}�� ���LC[ 42      W0���~��Q!��]�r��\      ��s���i�6 �eQ��      m�w�����Rv�=�      W~����!0Rf��C�h'      /s�n��<*����2iC!1      >kﳵ�i��*� ��h      y����u؎΂K (M�      wܮ����2�n
�      �:���1(��4I���Y[      ������� �/�?no      ��n�?��q��IȐj�      ������*`�)���){      /�=����d7�o%!      ���g703D
I�I�D      y��K�^J�7�5؁H�K      ����o$�8�6�b      o>�>�`lP�F��N+      nn���/��CBLCpH8�      S��Sz�����){        /�=�����d7 �o%!        ���g7 03D
�I�I�D        y��K�^�J�7� 5؁H�K        ���� o$�8��6�b        o>�>��lP��F��N+        nn���/����CBL CpH8�        S��Sz� X�t�ǀ              X�t�ǀ    