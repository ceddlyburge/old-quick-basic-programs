�(�  d0 0 ���^��8-��p8+-���      ���3��A�`�A�s�      k������z ܜz ��      �?����� `���d      ���5?�@f�� }��؟      ]������PQ  ��)Q��      ?�����r�� �r����      ?m������� 
�Ǿ���      Y������ � W�`����      �ǿT �$�@���v���      ]o��� �����{��      f���  �C(���g����      ����*� H	�� �K���      z�_�UU�`�W���p����      ������ �������      Ro�������������      ���U�.D���.�����      }�د��� '��������      ��a?��I�����M�����      ������L����\�����   UUK��  ���  �7��     
��y��  �X��  �_��     �����
�h"��
�l/��
�   /����.�_���_�O��_�  _��7�]����������  ���:>������������  ���|�|+�U��+�U��+�U  ������_� ,�_� ,�_�   �����t?� �?� ��?�   ���?����������  �������A_��A_���A_  /������z�C/�z�k��z�  �� �������������  ?�� ����W�?��W�$���W�  ?�� �������������  �@ ����B�������  ?�� ������?����s�����  �  ׃���(����;�����  ?�  ;G���?�����������  �  ��Ǉ�aǇ��c�Ǉ��  ?�  6��������� ������  �  �Ǉ�� �Ǉ� �Ǉ��  ?�  �����	���� �����  �  oǇ����Ǉ�@��Ǉ��  ?�  N�χ�����������;  �  _Ǉ�ޠ�Ǉ�'��Ǉ�?  ?�  ��ϯ�����
����
  �  �Ǉ�@�Ǉ��G�Ǉ��  ?�  �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            