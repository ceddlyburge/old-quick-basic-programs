���  d   �  �  �  �        x           �  H      �    � ��� ��      �           �  T        x  x        x  x        �  �       A� �       c� C�       3 #       ;��3��      ��      ?����      ?����      ��      ;� 3�       3� #�       a� �       @�  T        x          x       0  0  0     0  0  0  0  0  0  0    0  0  0  �  �  �  � ��������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        