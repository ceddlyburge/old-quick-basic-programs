��  d0 0 O����m���������  �  ������P?����S�����  �  {����Z�?���������  �  ������@���-�����/  �  ������ ���+������  �  ������ ?���������  �  ������ ��� ������  �  ��������������  �  >���������������  �  ���������'������  _�   /G�����G����G���  ��  _������������  ��  B����������@������ �  ��Ǉ���������� ��  ���C����� ����$ ��  ��?C����?C���?C�_ ?��  �@^�?�@^����@^��� ���  ����������������  ������C���CW���   �.�� �/�` �/�x����   _�� _��4 _��4����  ���>/>���?�����?������  ���|\���������������  ��@�?���@����@������@  ���t�����(����(����  UP���UP�DUP��6���     ���  �s  ��s���     ��w�  ���-  ������P   UUA��UU�2UU��:���   �����m���������ղ      ��������� A�����A      ���/������"t�����t      UT ��J��� ������ɿ        }�7���� ������        ��^���������       *������P  ����-       U_���f�� �����      ���g��   ؉E�����W      ������ $��=nC      ~��k���2D�e�:E�e      }������y����}�      �w�y��n�O�N~�_�N�      ��}��G ��
E����KU      ������ [f{Y�      ������H ��x&@���      ������@� ^	9c�^9;      )�̷}��;H� ��{H�       �zKo�K���߭��      �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            