�;�x;d0 0 ��> FCh�߹�Ch�߹�      ������ !
E���
      _���;ޠ
�'�0���?      M���e��,�%��,�%�:      k�����Ԁ B��[�C      �w����4� �u��      ��^��� �N��3?      7�S�y���%����-��      �?=?�l`���p�a�����      ;s�}����G笘�g[      ջ_?g*D����:t�ȱ�      ���?�� 8�?s%���      �|����� X �X<      ��_���I� ?�i� �      ����>?	��$ɚE��      ��x���'�T�'�TS      �����C 	�k�mP��      �p{ʻl�% ��% �  x   ?��!D���� �8    �� �?       �?���� ~  ?�9�      �����?��� <  �      �?����}� ?�}��?      �}��?����   G�~      �����x � ���~ @      ��~���  ���      ������ � ����~      ����~�q�  �| >      ���  3��@����      �3���`�`?o��  ��      p�`?�����><���9      ���=� ���8���?      ���������� ���      ������������� �� ��w�_�a��`��^�`����� ����� J�% �JDe    � f�׽���C(�DϹg���   � ]o������Hu��{Glu      �ǿo��$�@��v�@�O      Y��߿~� �"L��`��\�      ?m�������`A�Ǿ�eI      ?�����r��v�r���~      ]�����PQ��)Q��      ���5?�@f�� }��؈      �?����� `���d      k������z ܜz ��      ���3��A�`�A�s�      ���^��8-��p8+-���      �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            