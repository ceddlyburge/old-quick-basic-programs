�;�Ȝd0 0 ����,6�<��     �=��o|�A��� 2,��     �s�/�����x�H@���     ����kg�ژ^��x�u ߼     ���^�h@I�ה�9��:װ     yɸ��4�[� AlD���     um��~�hu�(dz���     if~�_�#E���C6!��h     7e՝����2|^�ˀ\     ��۲ �zh�5�3@@��     {�u�,� �g0ҷL���     ����~x�T�Ġ��     W�Ʈ}��n�s�ش
�|     ���N���F�,{����     ��޵/aJ����p��     �z�g��QO�4���      ��O���o-	$5�*Tl<     ��/]�k5zF	��
���      =�N����ie�Y `P0T�      �yu�c�q��!�@��a�l      ���5��ŷ(C4/�|�Ӵ      o�}�{�� 5�� ͼ      t�5?���d��`x�P�p      z�f�t��ֲ����ԛ�      <������1�a&�:
.�@     ?1�k?��B�	 H�      	R=Y���%�- B�fm��     �g���|�5l⑆z�`��     ��l-����h@hd�yp     _~����CMW�!���U      C�����:�L5�>��     M��}�=�7�� �{���      ���=���1�t�N��      �9���	��b�]      'k��=�5:@� j��À      �����y;@���]�����      ��z�m&	B�h���i��      [���n���*�߶�z      o׷�?w�)X����_NǛ      ��w��j������O�      �q߿��%�(r �'��z��      ٞsΐ�c�ޱ������      ���V�Va������_�      ~��3����̢�����      ڬ�~��'�� ��ᅳ�      O�|����T�r���|����      <�����Ӹ9)�ۿ�i�      Y�ݯ�<�{3]���{���      �o ��"JB        ���z�o `f�4 ���d��       �l����0n	i k��ʖ        ��2��� �8IXq m�*�        �}�z}� ��
��	 ���V        ��뽼_ %H�������"qh�       ��ئ�����.$�       �       ��.$��H(r��^|r��O�       ^|r��O�    