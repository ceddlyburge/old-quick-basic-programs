�;�p�d0 0 ����ym	$*��߮z�      �}�����Q� h_�Q���      �?����D�8F \���y      ������& !�Xawg����      ����͊A+c]2��;g��      �6���q�5X����O      �����Ch��g�;~�      ~__��v���p�����s��      ���~��H�1�xM�}      ��߼�ym0�����ώ�      5o���gް�L����      �����S	 �Ġ�몠     Ʈ޾�n�s�A��
�K�      ������FE3 {����      �޵���J�.�pn�     z����QO����@     ��O���o-	��*T9�      �/]�O�zFU��
�U��     =�N�o��ie�^ P0T�^      $yu�����!0B,�a>K�     }��5�=ŷ(t�/�|���      o�}�O}� 5��� ��      t�5�-Z�d�T�x�P��      z�f�o� ֲ��H����X      ������81�a�@�:
�R      �1�k��AB$!i H�j     iR=Y?^�%���2�f��      ��g���5l��z�`��      ���l��E�� �@hd��     �_~��n�CMW4����<�     �C����l�d@�L5���     �M����	�7�!1�{���     ��������1-��N=`     ��_}Y%	ű��Bb��     �gk����T5:A�j��0     �������)(@P��-h     ]ݟ���#�6+ &� ?      >��6��Qkia����q�     �������_���� ���     ݞ���"�mY� լO�     ����G�8SWx��R((���     z{����0�o�&"JB��     �z�o�~�4��d��     ��l���0n	iP�ʖ�X     2���_�IXq��*ħ�     �z}���
��	`��Vv�     뽼_�mH���ؐ"qh��     ئ���o�.$��    <�     �.$��o ��"JB        ���z�o `f�4 ���d��       �l����0n	i k��ʖ        ��2��� �8IXq m�*�        �}�z}� ��
��	 ���V        ��뽼_ %H�������"qh�       ��ئ�����.$�       �       ��.$��H(r��^|r��O�       ^|r��O�    