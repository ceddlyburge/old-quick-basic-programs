��rp �        ���        ���       ���   �   �?�  �   ��  �   ��  #�    � �   s�    ��   s�    ��   {�    � �   ��   �    
� U��U  �U 
��ʪ  ���   �    {�    � �   s�    ��   s�    ��   #�    � �   �    ��   �    ��    �    �?�         ���         ���         ���   U    
��   ʪ     �   ��         �          {�          � �         s�          ��         s�          ��         #�          � �         �          ��         �          ��          �          �?�                     ���                     ���                     ���                                                                                                                       