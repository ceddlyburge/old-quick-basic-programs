�;��@d0 0 ��2FCh� 9�Ch� 9�    ���^� �
E� a
  � _��";ޠj�'�0� F?  j� M��be��,�j��,� :  j� k��B}�ԀN�B��@ C  N� �w�Jo��(F� �` �  N� ��S~m� �F�N� 3?  ~� 7�Y�y���Ħ��� v�  � �?;�l`�ˍ��a�� s�  �� ;s�>:��
�G笀 g[  �  ջ+^g*D�ɐ�:t� ��  ;�  ���\�� I?s%� �  :]  �|vx���OX �  X<  v  ��i���IL ?�i   �  �l  ����>?q���$� ��  ��  ��,��� s�T� TS ��  ����C���k�  �� ��  �w4�}��Q`�� `� �X  ?�$3�wWY� ٜ ?.p  ﷿� �r@   ���  ��%��| x�@�   �����  {bj���xa�     �{c�  ������LT�   U����  ���}� Ά!   �e���   �g�����1A    1[��  ��|�����<J%   Z-+��|   ���� �JP   Z���   ����z�@@�  Aş��   �����~�B  ʺ���    p�x� �I�  i�� �    ��?������`  �����    �����   64��     >�� ��� ����>     ������ �"�"      z�_�f��`�R�^�p�[��      ����|� J�% �JE�e      f�׼���C(ÄϹg�ӌ�      ]o������Hu��{Glu      �ǿo��$�@��v�@�O      Y��߿~� �"L��`��\�      ?m�������`A�Ǿ�eI      ?�����r��v�r���~      ]�����PQ��)Q��      ���5?�@f�� }��؈      �?����� `���d      k������z ܜz ��      ���3��A�`�A�s�      ���^��8-��p8+-���      �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            