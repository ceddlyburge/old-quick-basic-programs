��rQ�        ���        ���     `  ���`   >    ���    >    ���    > p  ��p   >   ���    =�  �1    =�  ��    *� J��{   �z*��*�  x�� � � x�� � � �z*��*�   *� J��{    =�  ��    =�  �1    >   ���    >    ��    >    ���    >    ���        ���        ���         ���   �    �   �     �   ^�8   !T�   �T     �   !T    R�    ޫ�         w�     @    �C�         s�     @    �@�         x|          ���          |          ���          |          ���          |          ���          x          ���          8          ���                     ���                                                                                                                       