���  d              �   8  8  ?� :�   � p �    � p �      �         � @     � � 0  0  1� 1� `  `  a� a�       ��       �0�      �`�       ���@      ��ΐ      ����      ����      ����      ���@      �`�       �0�      �@        �  @ @  @  @� @  %@ '� '� '� 4  >0 >0 >0 ����     	        >  >  >  >                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         