���  d0 0 ^k��h}��ԟ������      �k���z�@D�nz�@��n      ���㿠<@�>1>l      |�߷���t`H*�~`ʪ�      �
��� 8( A08� C      @ ~�  �     `                                     "                   T T                   ����E                  UUQUU*                  ������                  _��_��                  ������                  ������            ��*��������            UUUUUU������            ������������            ������������            ������������            ������������            UU��UuUU��Uu�� *��      ������������UUUUUU      PUP UPUP U������                  ������                  ������      �    ��    �W����U      UU@UWUU@UW������      ꪐ
��ꪐ
��Uo�U       ��(����(�� ��        ���+�����+�� k�        ��DG����DG��  ��        ���/�����/��  W�        UW�_�@���_��  +�        *�꿮������  @        U�U �����  �         
��� ������  @         t}@ _����  �         ��� ������  @         |]  U��_�U  �          ��  �����  @          |\  ��_�   �        � �� ���  @       � |\  ��_�  �       � �� o���8 @       � || 0_��	8 �       ~ �� �/���� @       ^ || �_��� �       �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            