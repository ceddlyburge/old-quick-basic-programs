��r�K�        ���         ���    �`��`   �  ��#    <  ����    �p D��Gp   t  ����    � ��    � ��         ���         ���         ���         ���   3  D �D�   U"�"�   f  ��   u  ��   s  �   g  ��   U "�"�   6  A �A�         ���         ���         ���                                                                                                                                                                                                                                                                                                                                                                                                                 