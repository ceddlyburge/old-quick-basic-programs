�;���d0 0 �� d�2Ah� 9�Ah� 9�  d� ���$��  !
E� a
  $� _��$�ޠ"�'�0� F?  	&� M��4���,�2��,� :  6� k��4��Ԁ	��B��@ C  �� �w�0����� �@ �  �� ��_1�� ���N� ?  �� 7�1�������� �  �� �?9_l`؊�0�a�� 3�  
�@ ;s�9z���笀 '[  �@ ջFig*D���:t� 1�  �@ ���i{� #?s%� 6  k@ �|�Iw��1 �  <  y@ ��I_��I  ?�i   �  i@ ����^?	��$ɀ �  �@ ���O����  S  �@ �����C ��k�  �  �� �w٭}� � ���  �  Y�  ?�I�'w���®� �  M�  �+�$?��π�� �  _� ���$?�,BL��,S     Wl��|ߑ$<�"L� �f�     l�7�80��HL�>���    <L�>7�� ��ȁ��h@     <̡����N���E      Ώǿ��B h"��l+      J��y�rB��X�	���\�     K��K���1�� �|�2�     �1�����0 L�A�1�\�@     �1̶���cI�)� M�      �c}�.��� ͡� �     ������y.E�~.�      �Ro����푅�}����     /������L@� ���    /_��z�oLc��`��p�    /_k�����f: Q�% �@  %  �n f��N��CϹg�  �  _ ]o�L
����u��@  u  � ��L��$��v�v� O  �~ Y��@~� �L��`�  �  Y\ ?t�;������A�ǀ I  }ϸ ?���2��r���v�r� ~  }̰ ]���3�P!����  �  5ܰ �۔�/�@f1�� }� �  5�� ��o�����   =�� k�D[���	aܜ  �  e@ ���D_�A	a �A  �  e@ ��� -�8#p8+  ;�  #  �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            