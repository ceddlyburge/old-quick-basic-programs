���  d0 0 Hbٌ�=��9�³�����  �  �{���P�<߀ P����@  �  {�ٌ���"9��c���]  �  ����{�@X<ǔM\�����  �  ��ѭ�B�9��+�����/  �  ����~�<ǁ�-����  �  ���k?�XHk� ���k�  �  o���?�d<���o���s  �  6��c|��>c����c��  �  �]��nܘ�<ב'������  �  ���o}��	>o�T���o�\  �  3�Ƕw� ?����o����   �  ���m?�o� <�o��  �  �������� �����  �  �|�kA��>k� ;��k��  �  ���¨ *<����*����  �  ���i�@@i��a�i��  �  ������Q���Q����  �P ���X~�>X9��X  �����.���.���C�.��  ��T���T	�T���T  �����K�� �?K�� ��K��   �������W�*�W����W�   /��{��h
��a�
��c�
�   ���s�������ڌ?��   U�/_�_� ФQ�� Դ_��     
��߯-_�
 P�����_���     U^���롈 ���ȇ���      翿��E@@??�]S���      �m�� �� �������      ��_��� �  5����      ������ `  � ��,l��      ?�x��O�	�%���+�}ɿ      �����7D@/ �D@/�      �f���^z�J��{�ڟ�      _>����٠R  �٢R-       ��=��f�!��1˵�      Y�?g����؉E�6���W      o������I$��=nC      ~��k���2D�e�:E�e      }������y����}�      �w�y��n�O�N~�_�N�      ��}��G ��
E����KU      ������ [f{Y�      ������H ��x&@���      ������@� ^	9c�^9;      )�̷}��;H� ��{H�       �zKo�K���߭��      �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            