���  d0 0 ^ || �_��� �       ~ �� �/���� @       � || 0_��	8 �       � �� o���8 @       � |\  ��_�  �       � �� ���  @         |\  ��_�   �          ��  �����  @         |]  U��_�U  �         ��� ������  @         t}@ _����  �         
��� ������  @        U�U �����  �        *�꿮������  @        UW�_�T���_��  +�        ���/�����/��  W�        ��DG����DG��  ��        ���+�����+�� k�        ��(����(�� ��        ꪐ
��ꪐ
��Uo�U       UU@UUUU@UU������      �    ��    �W����U                  ������                  ������      PUP UPUP U������      ������������UUUUUU      UU��UUU��U�� *��      ������������            ������������            ������������            ������������            UUUUUT������            ��*��������                  ������                  ������                  _��_��                  ������                  UUQUU(                  ����D                  T T                     "                                   @ ~�  �     `       �
��� 8( A08� C      |�߷���t`H*�~`ʪ�      ���㿠<@�>1>l      �k���z�@D�nz�@��n      ^k��h}��ԟ������      �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            