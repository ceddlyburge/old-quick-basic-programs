���  d  � � � � � � � � ��������      � �     0 � �     0 � �       � �       � �        �  �        `  ` � � �    � � �    � � �      �  �   �  �   �  �        �  �        �  �        �  �    � �    � �    � � � �    �  �  �     �    @  C� C�    `  � �    0  < <    ���   ���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    