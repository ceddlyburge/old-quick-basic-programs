�;�@+d0 0 ��> FCh�߹�Ch�߹�      ������ !
E���
      _���;ޠ
�'�0���?      M���e��,�%��,�%�:      k�����Ԁ B��[�C      �w����4� �u��      ��^��� �N��3?      7�S�y���%����-��      �?=?�l`���p�a�����      ;s�}����G笘�g[      ջ_?g*D����:t�ȱ�      ���?�� 8�?s%���      �|����� X �X<      ��_���I� ?�i� �      ����>?	��$ɚE��      ��x���'�T�'�TS      �����C 	�k�mP��      �w�ʿ}�!5`���5`�      ?�v��w�Y�®��ٜ      �+�_���D@��   @  �����,B:B@�,S>��   @  |�����" E �f�    @  7������X@T����U�   �  7���}��`�!�h@ �e  �  ������D1AE  1[  �  ������h"�%l+ -+  �  y�x����X��P�\� �  �  K���z����2� �  �  ����}�L�C�\�P :  �  ����x�I�&�OM�  o�  �  }�4�{�� �2`� � ,�  �  ���y�.E2.�  �  �  Ro³�푮3��� T�  �  ����w� �"� "  �  z�F�f��`��^�p� �  �  ���T|� BF% �@ e  V  f��V{��C*dϹg� �  
v  ]o�N7���tHu��` lu  ~  ���o��$���v� O  �  Y���?~� �L��`� \�  �  ?d������`A�Ǡ eI  �  ?���n��r�v�r� ~  �  ]��
{�P?��  �  ?  ���B?�@fgP }� X�  g  �&��������� d  � k{���hύܜ` O�  
� ����A���A  s�  
ɀ ���-�8 @Rp8+  {�  A  �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            