�j�  d0 0 ƺ��P9E'2��9E'2��      ~:޳�?�šl�ؙե|��      �Z��z^0�Q��8��Q��      ���o�� �H:5�ȝ      �?�w���m�%�}�      ����_� 9� '���      k������0@@ �2O�G�      ����@������      ����3���*3����      ������
AU���      o>�_� ���������      ���'�  /��(<����      z���U�_�/������      �߄���W �_�_7����      ��KAEп��������      ��'�
�@!����@�����      |�_��������?����      �����������������      ���������?����    U��s�� ��� ?���    ������ i/��� i����    /����_���_����_��  ?�V���/B�(�/B�(��/B�  ?п�u���������?���  ?��{��	���	��?�	�  �����7���7��?�7�  ����<�P/���P/���P/�  ���}�w��Ђ���І����  ����������������  ���o�]��B�!���B�/���B  ���]���� ����'���  ���/6�����~�������  ���N�W�/� �W�/�#�W�/  �������^  ?�_a��_   ���?ۧ  =�,_  ?�=�  ?   ���i���~�?��=��   ��o�����"���"���   T ������)/���-����      ���_��(���;<����      ?;�
������������      ��  �!����%���      /�� ?�����ҿ���      [��UU}����6?���      �Ͽ���0@  62����      |������2   �2���      ����ϠP  8�5_��9      �k���z�@D�nz�@��n      ^k��h}��ԟ������      �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            