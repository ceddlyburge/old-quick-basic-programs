��r�        ���    8   ���   x   ���   |   ���   |   ���   |   ���  x|    ���   s�  @ �@�   w�  @ �C�   !T R� ޫ�   ^�8!T��T  �� ��  �� ��  �^�8!T��T  �!T R� ޫ�   w�  @ �C�   s�  @ �@�   x|    ���    |    ���    |    ���    |    ���    x    ���    8    ���         ���   �    �   �     �   ^�8   !T�   �T     �   !T    R�    ޫ�         w�     @    �C�         s�     @    �@�         x|          ���          |          ���          |          ���          |          ���          x          ���          8          ���                     ���                                                                                                                       