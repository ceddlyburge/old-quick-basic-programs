�;���d0 0 Dt嶣��!HP      ����2x���5wby      �}���k�Ɓ���      ��{�Η�|���F:Ԥ K      _���������L/� <Q:�      ����~��  $�kH���P      鮼���ɚ ݭ8� �"b      �ͺ���:�H �=a      �˴�?{R�����      �����΀1���xe�      �����"6=4Q�YƆ��       {�����DM�i3 �[��D      ��_��wH���F*D�P      ��+��W��h7p9��Z      ���u?���s#GP�=�X      ����Z�E��%a�x@8      �}��=c
d��@���      S����q7����*      �����# �bH      -��'MC�r4��0(*      G�r<����8���Vg0�      ��~���y�ۀ�ր��>A      ������1@z�@&�g       qf�w��%�p2F E<f(      �e�v3n#�kY]H�P��      k��{����0N�C��      ^�_��5)�������$      �����D!~ф�g3	      ��g3�(J
a���c=m�      �Zk}��� ���LC[ 42      �0���~#�Q!����r��\      ��s���i�6 �eQ��      m�w��ǅ��Rv�=�      �~����!0Rf��C�h'      /s�n��<*����2iC!1      >kﳵ�i��*� ��h      y�����؎΂K (M�      �ܮ���B2��n
�      �:��1(��4����Y[      �����x� �/��?no      ��n�?�.�q���IȐj�      ������*`�)���){      /�=����d7�o%!      ���g703D
I�I�D      y��K�^J�7�5؁H�K      ����o$�8�6�b      o>�>��lP�F��N+      �n���/���CBLCpH8�      ���Sz�� $ B        L��H5k �^����            ��
=�v��޳��T��  �       t������<��%�/            $�A$�" ?�̿��� `           �@�r��7�vޟu�
          d��1 w7z�o� "            #xG'�i�v)�~    �        !�$�Z     