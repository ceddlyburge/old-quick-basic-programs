���  d0 0 �zKo�K���߭��      )�̷}��;H� ��{H�       ������@� ^	9c�^9;      ������H ��x&@���      ������ [f{Y�      ��}��G ��
E����KU      �w�y��n�O�N~�_�N�      }������y����}�      ~��k���2D�e�:E�e      o������I$��=nC      Y�?g����؉E�6���W      ��=��f�!��1˵�      _>����٠R  �٢R-       �f���^z�J��{�ڟ�      �����7D@/ �D@/�      ?�x��O�	�%���+�}ɿ      ������ `  � ��,l��      ��_��� �  5����      �m�� �� �������      翿��E@@??�]S���      ^���롈 ���ȇ���      �߯-_�
 P�����_���     U/_�_� ФQ�� Դ_��     
��s�������ڌ?��   U�{��h
��a�
��c�
�   ������W�*�W����W�   /�����K�� �?K�� ��K��   ������T	�T���T  �����.���.���C�.��  ��T���X~�>X9��X  �ꀾ�����Q���Q����  �P ���i�@@i��a�i��  �  ���¨ *<����*����  �  �|�kA��>k� ;��k��  �  �������� �����  �  ���m?�o� <�o��  �  3�Ƕw� ?����o����   �  ���o}��	>o�T���o�\  �  �]��nܘ�<ב'������  �  6��c|��>c����c��  �  o���?�d<���o���s  �  ���k?�XHk� ���k�  �  ����~�<ǁ�-����  �  ��ѭ�B�9��+�����/  �  ����{�@X<ǔM\�����  �  {�ٌ���"9��c���]  �  �{���P�<߀ P����@  �  Hbٌ�=��9�³�����  �  �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            