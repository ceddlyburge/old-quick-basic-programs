���  d0 0 P�/ �?�/�� �       ��^�	p_�_�p �       x�? �?�?� � �       p�^��_�_�� �       ��/@  ?�/�0 �       X�� �_���0 �        x�/@ �?�/� � �        t�� �_��P� �        8�/@ �?�/��� �        ��� _���4 �        ��/�  ?�/��  �        d�� �_���� �        l�� �?���� �        8�� �_���� �        ���P(?���j �        L����_���� �        ,�
���?�
��� �        X���_��� ��       l~��������� }P       | �@U��/�@U��  ��       d~�
����
�� _�@      � �@U/�@U  ���      z � *��� *�  W��      ~ _�  ���  �  *��      t /� ��� �  _�      � �J (��J *  ��      � �������   U      � ��Uh	���Uj   �      ��������           �� �������          @ U_���������          }� ���A_����@          �`  UU@�����@�          ��  
� ���`          ��    W +���_�          z�    ������          ��     ����(�          o�    � W���          _�   �� )UUʮ          �5�   � ���          �(   ��   ���         k��   �(   �},         ��  BD   BN�        ���,  !H�  %!��        ���w���H:5�H�      �Z��z^0�Q��8��Q��      ~:޳�?�šl�ؙե|��      ƺ��P9E'2��9E'2��      �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            