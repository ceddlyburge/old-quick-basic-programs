���  d  � � � � � � � � ��������       �  �     `  �  �     `  �  �       � �        �  �        x  x        0  0  �  �  �    � � �    � � �    � � �  8 ������ 8 ������ 8       8  8       � �       � � ��� ��� �    � � �    � � �@  @�@ x  x�  � x�     @ � �     @ � �     � x� x�   ������   �@�@�@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    