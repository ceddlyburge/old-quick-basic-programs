�D�  d0 0 ƺ��P9E'2��9E'2��      ~:޳�?�šl�ؙե|��      �Z��z^0�Q��8��Q��      ���o��  �H?���ȝ      ����w�   m����}�      ����_�   9� ������      ������  @ ����G�      �����UYP�������      � �����*������         ������AU�����       U _� �����������      U��'� �����������      ����U����/�������      ���������_�������T    �_AE�_����_���k��   @ /�
�@ /���@ /������   �T���T����T���o��   +�����+�����+��������   _�E���_�E���_�E������ U����� ����� ����� ��� ����� ���� ���� ��� /��W�_���W�_���W�_������V��/B���/B���/B����п�������������������@�	��@�	��@�	�������P���7�P���7�P���7��_����qP/�qP/�qP/�����������������������[�?��[�?��[�?���������W��B��W��B��W��B ������5����5����5�� ������ ���� ���� �� ����U] W�/�� W�/�� W�/ ���Ъ���^����_����_ W�����  =���  ?���  ?  	���P�`~���`���`  ����_���J�����������   UT ��+��� ����������      �`_�� �����������      �� 
� U����������      �   � ����������      ��� ?� U��������      [��UU}�  ���7�����      �O�����   6�����      |������p   �����      ����Ϡ  8�>?��9      �k���z�@D�z�@���      ^k��h}��ԟ������      �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            