��6 d0 0 %�m�$�
���      ���� O3A�Fx��      �wx� �c�@ i���      �s��� /�k>���%+W      ��o?� �2��q\�<,      �~�?� �;$��
9zs      �;'=` �� Y�FDm-�      ��m]� \@�-�t��M +      ���-� cE�I0Sٶ�      sWM�� ������K      �����@Y�,�lD�ac�      ]���o�̖�"�"e���       ��������=��
G"Tb�      ��?�㓜�+A`�Z7��      ���7��@����3�i
�      Z�������a�S��      Ƽ��S�&P�Ȁ���      ���У�!i�@�T�� 8      u���`��ĽX��F !      ���x1��M,N��T`       �]<N�����Q�jA�      Y��~��)�E�@�|/�k      �}��k�X^� @�Ad      �X�_f�bL����f<�      v�n��������W
s@      ���{���8�H���Cr      ����zp���$-      5x�-��H�~�"��昃!      �����#mY�PR���+      m���Z?2��EiL,��      ~�����e����:+N��      �o����@� l���Xe��      ��e� ��#�[nJ      ���{~�fJ��0��p      �1v���G!I5T<@��L      G����|�XT'�����      ���畞�Asq�W� �      ��wu;��LBPv��      ����\�,A�� ښ�3�      �ۿ����c ���v�A      ���v�_5m��3tkV	��      ����=Ք9T�((�Q�      ����W��&w��������      �����X`P"�"M�A'�      zm�c�- ��Rҧ��      �������5$8�Fp��l@      �|��|� 
�6�rqbp      �{{�vw2B�%QI-��      ?^�7_�� $ B        L��H5k �^����            ��
=�v��޳��T��  �       t������<��%�/            $�A$�" ?�̿��� `           �@�r��7�vޟu�
          d��1 w7z�o� "            #xG'�i�v)�~    �        !�$�Z     