���  d              �   8  8  ?� :�   � p �    � p �      �         � @     � � 0  0  1� 1� `  `  a� a�       ��      �0�       �`�@      ��Π      ���`      ���@      ���@      ���`      ��Π      �`�@      �0� @  @  C�AH`  `  `� `@  �  �  �  � *P@?�@?�@?�@5�?��?��?�� 
� � � �0�0�0�0� � � � �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                