��r�0�        ���        ���       ���       ���       ���       ���        ���         ���      ��� O      ���     0 u�8�    y����    K0{�>�    y����     0 u�8�       ���       ��� O         ���         ���         ���         ���         ���         ���         ���   K0   {�>����          y�   ������           0    u�8����                ������                ������ O                  ������                  ������                  ������                  ������                  ������                  ������                  ������               ������                  ������                  ������                  ������                  ������  