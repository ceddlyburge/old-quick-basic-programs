�;�8�d0 0 _�!P�D!   �@     !P�����qwbyu     ���s�k�Ɓ�1��0     {�Η/�|����Ԥ K�P     ����w��L/Ȁ<Q:�Ȁ     ��~��� $�k��PX      ����ٚ ݭ& �"b4�      :���wzt:����=aϭ�     �?{]����Ʋ��      ���U����/xe��.     ������=4Q� "���  �      ���j?̀i3��[��D��      _��wG1����*D�P��      +��W]�h7p9�A�Z�@     �u?-��s#��=�X�X     ��Z;m��%a̐@8ΐ     ��=c�
d�������     �����q7�����*�     ����w��#�bH�     �'M��r4��:60(*:0     r<��}�8���*Vg0��(     ~���1��ۀ�� ��>A�     ������z� 2�g (0     �w�=ݭp2F�!<f(�      �v3n{5kY]���P����     �{��\��0�\C����     _��5~�����贈$��     ���w�~ъVg3	�V      g3���
a��c=m��      k}��(�⏋L� 42ד      ;��~��Q!��9 ���\9!�     3���[�� ��KQ�ť_      w���~����=���      ������Rf��`�h'`      �n��{�����C!1�      o���]��*��@��h�@      '�����΂K[ (M�[�      �����|��n
��      ����(��40���Y[0�     ���l] �/���no��     n�?�u�q����Ȑj֋�     �������)��x@){xL      �=��m�d7��%!��     ��g7OD
�I�D��     �K�^{m7����H�K�     ���:,$�8����b��     �>�v|P�����N+��     ���/?�CBL�0H8��     �Sz��� �B){�xH      �=���m�d7 ��%!���      ��g7�O{D
��I�D ��      �K�^�{m7� ���H�K�m�      ����:,$�8� ���b�U�      �>�v|P� ����N+���      ���/�?�CBL��0H8� �      �Sz����e�  a�w         �����    