�j�  d0 0 �Ǉ�@�Ǉ��G�Ǉ��  ?�  ��ϯ�����
����
  �  _Ǉ�ޠ�Ǉ�'��Ǉ�?  ?�  N�χ�����������;  �  oǇ����Ǉ�@��Ǉ��  ?�  �����	���� �����  �  �Ǉ�� �Ǉ� �Ǉ��  ?�  6���������������  �  ��Ǉ�|aǇ��c�Ǉ��  ?�  ;G���8�����������  �  ׃��� (����;�����  ?�  ������?����s�����  �  ����B�������  ?�� �������������  �@ ����W�?��W�$���W�  ?�� �������������  ?�� ���z�C/�z�k��z�  �� ����A_��A_���A_  /���?����������  �����t?� �?� ��?�   ������_� ,�_� ,�_�   ���|�|+�U��+�U��+�U  ���:>������������  ���7�]����������  �����.�_���_�O��_�  _�����
�h"��
�l/��
�   /��y��  �X��  �_��     ��K��  ���  �7��     
��������L����\�����   UU��a?��I�����M�����      }�د��� '��������      ���U�.D���.�����      Ro� *�����������      ����   �������      z�_�  �`�W���p����      ����T  H
�� �K���      f������C( U�g����      ]o������   ��{��      �ǿ��$�@� �v�@��      Y��߿~� �"L��`��\�      ?m�������`A�Ǿ�eI      ?�����r��v�r���~      ]�����PQ��)Q��      ���5?�@f�� }��؈      �?����� `���d      k������z ܜz ��      ���3��A�`�A�s�      ���^��8-��p8+-���      �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            