�;�(�d0 0 �� d�2Ah� 9�Ah� 9�  d� ���$��  !
E� a
  $� _��$�ޠ"�'�0� F?  	&� M��4���,�2��,� :  6� k��4��Ԁ	��B��@ C  �� �w�0����� �@ �  �� ��_1�� ���N� ?  �� 7�1�������� �  �� �?9_l`؊�0�a�� 3�  
�@ ;s�9z���笀 '[  �@ ջFig*D���:t� 1�  �@ ���i[� #?s%�   k@ �|�Ig��1 �  <  y` ��Ig��I `?�i   �  i` ����6?	���$ɀ �  �� ��̳���P�   S  �� ���͙C �x�k�   �  �� �w٭�}� �<���  �  Y�� ?�I�fw��®�    M�~ �+�%��ώv��     _�v���$��,BLǿ,S      Wl��|ߑ$x?�"L� �f�     l�?7����HL�����     <L��7����Ȝ��h@     <������O����E      Ϸ����B�h"�l+      J�y�rB8��X�	���\�     K��K���x�� �`�2�     ������|�L�A�?\�@ 0   ������pwI�)�FM�  `   �}�.�y�� ͡� � (   ������x�.E��.�     � �Ro����푅���� T�  /�����L�� �"� "  /^� z�oLf��`�^�p� �  /_@ ����|� Q�% �@ e  �@ f��N{��CϹg� �  _@ ]o�Lw����u��@ ,u  �@ ��Lo��$���v� O  �@ Y��@~� ���`� �  Y` ?t�?������A�ǀ I  }Ϡ ?���.��r���v�r� ~  }̠ ]���;�P!����  �  5܀ �۔�?�@f1�� }� �  5�� �������   =� k�D;���	aܜ  �  e  ���D�A	a �A  3�  e  ��� -�8#Rp8+  {�  #  �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            