�;��qd0 0 _�!P�D!   �@     !P�����qwbyu     ���s�k�Ɓ�1��0     {�Η/�|����Ԥ K�P     ����w��L/Ȁ<Q:�Ȁ     ��~��� $�k��PX      ����ٚ�ݭ& 6"b4�      :���wzt�:���2=aϭ�     �?{]����Ʋ��      ���U����/xe��.     ������4Q� "ę�  �      ���j?πi3��ݍ�D��      ߍ�wG1���ϮD�P��     ���W]�x7p9�C�Z�@     �u?-��s#���X�P     ���Z;K��%a̜N8΀     ��=c)t������      9����x�w��{�*     {����C��#��"H�     ��'M<v4��qð*      }��<��?�����0�      ���������ۀ�<8�t>A      �����������g       ��w���p2F��f(      ��v3n��kY]��P��      ���{��`<�0>~��      >~?��5p0��p00$      p0?��<8b�  }g3	      <8g3��8!��?�m�      ��?��� ��Lp7� 42      p7���~?��ᦫ�� �\      ?�����q0 �r ��      s0��� ���z=�      �~����9��A��'@     ?�y�����1�     �����\
l*�����h�      �����>΂K[(M�[�     >����v��n
��     ����+��40��XY[0�     ���lY �/���no��     n�?�u��q������j֋�     �������)��x@�{xL     �=��m�d7���%!��     ��g7O@
��I�D��     �K�^{mX7����H�K�     ���:,d�8����b��     �>�v|P�����N+��     ���/?�CBL�0H8��     �Sz��� �B){�xH      �=���m�d7 ��%!���      ��g7�O{D
��I�D ��      �K�^�{m7� ���H�K�m�      ����:,$�8� ���b�U�      �>�v|P� ����N+���      ���/�?�CBL��0H8� �      �Sz����e�  a�w         �����    