�;�`�d0 0 �!HP	@t!         �!HP	�x���(5wby      �}����k�Ɓ��      ��{�Η�|���F:Ԥ K      _���������L/� <Q:�      ����~�)  $�kH���P      i���� ɚ ݭ8� �"b      8ͺ���:�H �=a      �˴�?{�R����n���      �����΀1���xe�      �����"6=4Q�YƆ��       {����[DM�i3 �[��D      [�_��w���F*D�P      ��+��W��h7p9��Z      ���u?(��s#GP�=�X      o���Z�E��%a�x@8      �}��=c
d��@���      S����q7����*      �����# �bH      -��'MC�r4��0(*      G�r<��1�8���Vg0�      3�~����y�ۀ�V���>A      ������1@z�@&�g       qf�w�e%�p2F E<f(      ee�v3n#�kY]H�P��      k��{����0N�C��      ^�_��5�)���0���$      ������!~��g3	      ��g3٨J
a��Tc=m�      �Zk}�� ���LC[ 42      W0���~��Q!��]�r��\     ��s���i�� �e��     m�7���}���Rb=� `   W ��&��f��	"h	�� �(  n�0����/ c� oP    ������   �  @      �>�m�3d��L�~ɗ���      �:����(�{�
?���
      �|������k����v      ���_�	���뵤      ���~��)�� ti���L      ^<~����ÃU� ���׺�      �U�_�.,��P�m�n���      =^��¡6X�v�?>~�      =�?�]o�M�&�Wm����      �xs���+��s[?����[      ������B�fo^M�E�      ������)+�7mo�_�      ����ÃU�  ���׺��       wU�_�.����P� m�n��� �      =^���¡6X� v�?>~��       =�?�]o��M�&� Wm�����       ]xs�������s[ ?����[ �      }����݀��f o^M�E� �      �������)+� 7mo�_�        ������       7�sN���           