�;���d0 0 �!HN�@t!     �!H@ �x���(5wh*    n�}�� �k���C    珋{�� �|���F:ԤP    �_���� ����}�� <Q�    �����@ )  $��H���a    vqi���  ɚ ��8� ��    O�8ͺ�  ������H �l    |��˴�  �R��}�n���A    �G����  �1��]��x��    �����  "6=4��YƆ�,    l�{���  [DM�] �[���    >�[�_�� ���_�F*D�,    s,��+�� ��h7_��Z �     ����@ (��s7wGP�=Ȩ    �o��� �E��;�x@L    ��}��  
d�}@����    �S��� q7�;�� �    ���� �=� �bD    t-��  C�r4��0(!    %G�r<� 1�8����Vg/    �3�~�� �y�۟�V���     ����� 1@z�@&�g    �qf�w  e%�p7� E<f    ee�v  #�k}�H�P�    {k��{� ��N�C���    �^�_�� �)���0���     X����  �!~w��g     ��g  �J
a��Tc=      D�Zk}�  ����C[ k     k�W0��  ��Q!��]�r� i    �k��s�  i�6��eQ�$   mm�w�  ѻ�Rv�<D$   �wW~��  !0Rf��C�iS   �/s�n  <*��92iC Ƅ    ��>k�  i��*�� �J     �y���  u؎η (L�    �wܮ�  �2��n$    6�:  �1(��I����    +������ �� �_|?n �    (���n�  ��q�IȐ.�    ?ܿ��� *`�)���)	�    �/�=� ����o%     5���@ 03D
?�I�I��    �y��K� J�7�5؁H�*    {��� o$�;�6�    o>�  `lPקF��HX    �nn��� ��C^�CpH!H    �S��S` �߀�)	�     � /�=�  ��߀�o%      5 ���`  03D
��I�I��     � y��K�  J�7��5؁H�*     { ���  o$�;��6�      o>�   �lPק�F��HX     � nn���  ���C^��CpH!H     � S��S`  [ON���              [ON�      