�j�  d0 0 �
�]c7�L䢜7�L䢜      ���{\~6���;e>���      z^w�Z󕡊�����      _�����	 (�H�\      ��O��_���7�闤      ��c��� ��0������      ������ �)����L�      W������ !��/�0i      ����{�T!!�0�����0      U�/������P�����S       ��|��@�	�����       W������0����<      ���^��/��������      U�!������������      �����?����������      �P�{�����������      ����>����@�������      ���_������������      U��/U����U���઀     ?��� ?���  ?���8�� 0   ���i ���� ������ x  ��������������j�  �B����B���B�����  ��X���X�Q��X������  ���?�����!����w��_�  ��G����G���G����  W�
�<wW�
�ÈW�
�������  �W�W��A�W��a����  ����?���������������  B��{�B����B��������  ���8�����?E���?�E_���  ��ul���~����ߋ���  �/�p�r�/���/�ď���  z@����@� �@�����   �  ����  �4��  �����   ~�������(i�����_�   ��W����W�D	��W�D *�   ���K{���ؔ����ش      �_���'?��������<�      �-P�����#�����[      �  /���Є�?�����      � _������K�����K�      ������AUU@�%o����l      �����  @����Ll      _����>�   L�����L�      ����_�  
��_���E      ����ֿvW"-^vW��^      ���zA�+�/�E�����      �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            