�;�Qd0 0 ��0��Ch�!9�Ch� 9�  �� ������ 1!
E� !
  �� _����ޠ5�'�0� ?  �� M����,�4��,� :  �� k�����Ԁ�B��@ C  �� �w͒���1� �p �  �� ��]E� ��rN� ?  �p 7�Qa����z��� �  �x �?<��l`��w��a�� �   �� ;s��:�笘 [   �� ջ^��g*D�3��:t�  �   �� ���x�� 80�s%�     x���|��W����  <   _���I�`�I���i�    �`����c�	f0$ɚ@    g���v<��'׿�'�    ������C 	��k�mP     ���p{ɣ�!B`�     x�l?��1��   �   �81�  �� �?       �?���� ~  ?�9�      �����?��� <  �      �?����}� ?�}��?      �}��?����   G�~      �����x � ���~ @      ��~���  ���      ������ � ����~      ����~�q�  �| >      ���  3��@����      �3���`�`?o��  ��      p�`?�����><���9      ���=� ���8���?      ���������� ���      ������������� �� ��w�_�a��`��^�`����� ����� J�% �JDe    � f�׽���C(�DϹg���   � ]o������Hu��{Glu      �ǿo��$�@��v�@�O      Y��߿~� �"L��`��\�      ?m�������`A�Ǿ�eI      ?�����r��v�r���~      ]�����PQ��)Q��      ���5?�@f�� }��؈      �?����� `���d      k������z ܜz ��      ���3��A�`�A�s�      ���^��8-��p8+-���      �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            