�;� �d0 0 Dt嶣��!HP      ����2x���5wby      �}���k�Ɓ���      ��{�Η�|���F:Ԥ K      _���������L/� <Q:�      ����~��  $�kH���P      鮼���ɚ ݭ8� �"b      �ͺ���:�H �=a      �˴�?{R�����      �����΀1���xe�      �����"6=4Q�YƆ��       {�����DM�i3 �[��D      ��_��wH���F*D�P      ��+��W��h7p9��Z      ���u?���s#GP�=�X      ����Z�E��%a�x@8      �}��=c
d��@���      S����q7����*      �����# �bH      -��'MC�r4��0(*      G�r<����8���Vg0�      ��~���y�ۀ�ր��>A      ������1@z�@&�g       qf�w��%�p2F E<f(      �e�v3n#�kY]H�P��      k��{����0N�C��      ^�_��5)�������$      �����D!~ф�g3	      ��g3�(J
a���c=m�      �Zk}��� ���LC[ 42      �0���~#�Q!����r��\      ��s���i�6 �eQ��      m�w��ǅ��Rv�=�      �~����!0Rf��C�h'      /s�n��<*����2iC!1      >kﳵ�i��*� ��     y��� �؎΃} (L�     ��ܮ�� B2�˕n
v    ��:� 1(�������P"    >����� x� �+?�?n�    ���n�0 .�q��IȐa    R����� *`�)���)    ,/�=� ��o��o%E    g���` 03D
�I�I�I    Ky��K� J�7�5؁H�	    ���� o$�;�6��    �o>�  �lP�+F��R�    ��n��� ���CG�CpH:     ����S` � $ B        L��H5k �^����            ��
=�v��޳��T��  �       t������<��%�/            $�A$�" ?�̿��� `           �@�r��7�vޟu�
          d��1 w7z�o� "            #xG'�i�v)�~    �        !�$�Z     