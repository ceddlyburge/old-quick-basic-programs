���  d0 0 ���^��8-��p8+-���      ���3��A�`�A�s�      k������z ܜz ��      �?����� `���d      ���5?�@f�� }��؈      ]�����PQ��)Q��      ?�����r��v�r���~      ?m�������`A�Ǿ�eI      Y��߿~� �"L��`��\�      �ǿo��$�@��v�@�O      ]o������Hu��{Glu      f�׼���C(ÄϹg�ӌ�      ����|� J�% �JE�e      z�_�f��`�R�^�p�[��      ������ �"�"      �o������������      ������  ��64�      ������  `�����       ��x��� I�������      �����������ʺ      ��Q��z��� ������      U�����U��
PU����      ��w�� ���% ���-+�P    �U-���U/�1A�U/�1[���   �P�}��P��!�P��e���   ��G�����T����U����   ң���� �� ���   �*�W���*�x@��*������  �t����t�@�t�*��@  ~�s�w��|Y���ٜW��  ��/'�}��/8`���/?`� 
��  ��W����x������  �   C#����C<T��C?TS  ��  ���s>?�|�������  /�  ��o��� O� ?��� �  @  ���W�� �xX ��X<  �  ��m�����?s����     վ�sg*A�|��:���  �  ;vk3����<G��?g[  �  �>�c�l`��|p�a����  ?�  7�c3����<&���?��  �  ������ ��O�߳?  /�  �~c3����< ��?��  �  k�����ԁ��B�����C  �  M�c3���)�<�/�?�:  �  _�1��ޠ�D'�7��?  �  ��[3�� �<!
G�?�
  �  ��1�FCh��Co��  �  �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            