��rh�        ���   ?@  ����  >� A ��  ]� " ��  k�  ��  t�  ��  o@ � ���   ?@  � ���         ���         �f         ���         ���         �w         �f         ���    �   ��    =�  ��#    � 0`�pc    '` ��؃    2` ��̓    <�  �C    �  �d         ���         ���                                                                                                                                                                                                                                                                                                                                                                                                                 