�;��d0 0 � B ����w:            X
����W�            �"�
,���}m�            b2����5�r            h�A �v�>�             0!B�����             $`H� �ە�             ~�����            `�B  �0�a�            "!(D  �V�;]�             Ar�]���             ЀP��n��            �8@�u�w��            ��$��}��v�            a!�זH���            �@��)���            � &@"o�"���            JA�@Y5���            @&�h �ةO�              � k�x�D�            !���z���              @� Ϸ�+S�            �B] �l���             QR]����i            ��  �}�w��            "�  ���[��            � �h�n��Y             	 �sb;,}�            �   $6ݱ��            ����~E�~            @` �;k��o             @ `�����u             �D��[؍#            ��
,L ~����            �PX ��l,���e            Hp @����ӽ            �  C��[۟��            ����y�_�m�              `��<�����            IP �r���_            @	`! @����            �@%Ѐ�t?�qo            � �"B��_Y�              @A0�ޏ���             A)@ B�/���             ��@�]��2              @!�!�ϟ�|�            $ I�hڻ��#                                                                                                                                                                                                                                            