��k6 d0 0 |�> F�h�߹��h�߹�      ������!
�U���
     ����;�` 
�'z2���? 0    �k��e�r�%�s��%�: �    k�v����� B��۬C r�   �7��
�� ����R�   {�~���� ����3?S@   ����y�
 %����-��U�   ^�-?�l���p��������   �_�}��$  �G/���g[ �p   _��?g�  ����}�ȱ�u�   o��?�̀  �?������>   p�;��߀  X ���X<�   ^��_�� � ?���� � ��   ?���>?� �����E��~    \x��� '�T����TSـ   x����� 	����P��|�   ��ʿ}G 5`�O��5`��8   o�~��w� �Y�ӿ��ٜ�   3����DD"@����    ��]���(@*"@�/{�.��)�   ������  o� (�   7�|�?��X�h�����h�      7����� �	�hE�U�     ������` Ez2�    0 ���k�h"r�l+s��    � y�k�w�X���
�\����    r�K���7~�
��2���   R����{�L�H� �\�Z���   S@������I�"
!M�"��   U�}�?^�-� Ѡ ����   �����_�.E $  .�6/��    �pRo�_��푤� ����}�   u����o�� �  ����   �>z�_p�;�`�� �p����   ����^�� J�  �J���    ��f��?���C(� �g����   ~ ]o�\��� '��{���   ـ��x�ր$�� 	�v����   |�Y���� �G �`�O��   �8?mo�~���� ��Ǿӿ�   �?��3��r�DD�r����   � ]����]�P(@*��)/{�   )�������@f }�o�   (��?����� `���d      k������z ܜz ��      ���3��A�`�A�s�      ���^��8-��p8+-���      �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            