��rX|�        ���        ���       ���       ���       ���   �   �?�   �    �?�    �    ��   `�    ��   0�    �?�   �    �?�   >��   �    >��   �    �    �?�   0�    �?�   `�    ��    �    ��    �    �?�    �    �?�         ���         ���         ���         ���         ���                                                                                                                                                                                                                                                                                                                                                                                                                 