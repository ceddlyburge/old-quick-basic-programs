�V�  d0 0       
��                     U�                     /��                   W��               
��   ���               W@   _��               ��   ���               ��   ?��              W�   �W�    �          ��   ~��   U          E�   �E�    �          ��   ~��   }          E�   �E�    �          ��   >��   U          u�   �u�    �          �@   ?��              ��   ���                   _��               ��   ���                U    W��                     *ݪ                     UT                     
��                     UP                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               