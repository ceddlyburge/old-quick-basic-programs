��r�%�        ���   �   �?�   �   ��   �   ��   x   ��   |   ��   >    ��   p?    ���   8    ���   , 
����   ���  ��  �   ��  �   ���  , 
����   8    ���   p?    ���    >    ��    |    ��    x    ��    �    ��    �    ��   �    �?�         ���   ��        �         ��      �        ,    
�   ���         8          ���         p?          ���          >          ��          |          ��          x          ��          �          ��          �          ��         �          �?�                     ���                                                                                                                       