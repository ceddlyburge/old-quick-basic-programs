���  d           � � � �  �  � ?� 
�  @ @ s� -@      q�        }� "@       ?�    @  @ � @  `  ` |` |`  0  0 �0 �0      A� A�       c� #�       3? ?       ;��+��      ��7��      ?����      ?����      ��7��      ;� +�       3? ?       a> !>     @�@�  0  0 x0 0 (  x  x  x R�����`������
� � � � 
 ` ` ` `                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        