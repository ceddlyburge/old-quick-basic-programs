�;�HFd0 0 ��&�Ch�	9�Ch� 9�  � ����� �!
E� a
  �� _��,�ޠD'�0� F?  -� M��l���,��,� :  m� k�����Ԁ�B��@ C  ɀ �w�<���,s �` �  � ��A�� �RN� 3?  V� 7�C0����r&��� v�  r� �?#0�l`��b0�a�� 3�  r� ;s�z���笐 '[  �@ ջT��g*D����:t� 1�  �� ��Ĕ�� 6ք?s%� 6  �� �|������� �  <  �� �蟿��I��?�i  �  �� �����?	���$ɘ �  �� ������!�d�  S  �� �����C 	cr�k�h �  �� �w�u�}� 1����  �   u� ?�t\�w�Y��®� �   ]� �+�nǀ�DL� ��      n����`s�,B:fs�,S>      fs�|��# o�" � �f�      �o7�1�8��Xp�����      q��7��w�� 0q��hE      1w������E      ������h". l+      �y����X�'��\�      7�K���� �A� �2�@     � ������L�H@?<\�Z�     �������I�"H�M�"h      ��}�?�@ � �? � �       �����.E  �.�64      �Ro�`푤�������      ������ �"�"      z�_�f��`�R�^�p�[��      ����|� J�% �JE�e      f�׼���C(ÄϹg�ӌ�      ]o������Hu��{Glu      �ǿo��$�@��v�@�O      Y��߿~� �"L��`��\�      ?m�������`A�Ǿ�eI      ?�����r��v�r���~      ]�����PQ��)Q��      ���5?�@f�� }��؈      �?����� `���d      k������z ܜz ��      ���3��A�`�A�s�      ���^��8-��p8+-���      �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            