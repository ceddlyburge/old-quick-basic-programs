��r���        ���    �p  ��p   �  ��   �p  ��p   �@  ��@   �p  ��p   �   ��    �   ��         ���         �fg         �ww         ���         ���         �fg         ���   �    ��   �    ��   �    �g   �    �w   �    ��   �    ��   �    �g         ���         ���                                                                                                                                                                                                                                                                                                                                                                                                                 