���  d0 0 ��1�FCh��Co��  �  ��[3�� �<!
G�?�
  �  _�1��ޠ�D'�7��?  �  M�c3���)�<�/�?�:  �  k�����ԁ��B�����C  �  �~c3����< ��?��  �  ������ ��O�߳?  /�  7�c3����<&���?��  �  �>�c�l`��|p�a����  ?�  ;vk3����<G��?g[  �  վ�sg*A�|��:���  �  ��m�����?s����     ���W�� �xX ��X<  �  ��o��� O� ?��� �  @  ���s>?�|�������  /�   C#����C<T��C?TS  ��  ��W����x������  �  ��/'�}��/8`���/?`� 
��  ~�s�w��|Y���ٜW��  �t����t�@�t�*��@  �*�W���*�x@��*������  ң���� �� ���   ��G�����T����U����   �P�}��P��!�P��e���   �U-���U/�1A�U/�1[���    ��w�� ���% ���-+�P    U�����U��
PU����     ��Q��z��� ������      �����������ʺ       ��x��� I�������      ������  `�����      ������  ��64�      �o������������      ������ �"�"      z�_�f��`�R�^�p�[��      ����|� J�% �JE�e      f�׼���C(ÄϹg�ӌ�      ]o������Hu��{Glu      �ǿo��$�@��v�@�O      Y��߿~� �"L��`��\�      ?m�������`A�Ǿ�eI      ?�����r��v�r���~      ]�����PQ��)Q��      ���5?�@f�� }��؈      �?����� `���d      k������z ܜz ��      ���3��A�`�A�s�      ���^��8-��p8+-���      �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            