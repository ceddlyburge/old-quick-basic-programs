���  d0 0 �
�]c7�L䢜7�L䢜      ���{\~6���;e>���      z^w�Z󕡊�����      ?�����ЀH(րL�\      ��{_� ���� ���      � k��@  �B0@ �B�         ���  S)  ���         ��� P?8!   ?;i         ;����$0   5S0         '��UW�%   eS         �����	   /         �����            �^����c�   
c�      uT�������   ��      *���?�����   ��      U��������    �      �����>�����    O�      ����������   	�      ����s������   ��      �UW����UW�*  �� j8      �����i����
�UUTJ�      U ��U ��������         �>�   ����� �         �_�   ��Q�����      � 
�Pު 
��!U�� �w      UUU���UUU������      �����w���� �UT (�      �����������A   �a      ����������    ��      ����?�������    ��      U��A}������E    �E      *����������   ��      UU�r����D�   M�         ,������   ۆ         ������!�   /�         �W��
�i   
��         ���UT	            /�{����   ʴ         =�'U@C�   s�         ��� *�B   NG[        ��   WE�   �e�        [��  �A�  �ˑ        �ڀ  �8%� "�8l      m���R��$�@�$�l      �����>@T.��US~�      ������<�(6|��|E      ����ֿvW"-^vW��^      ���zA�+�/�E�����      �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            