���  d0 0 � ��
@/��@ �       �z/@p_�/�p �       � �� /��0 �       �z/@@_�/�� �        ������ � �        x/@_�/�  �        �����  �        �/@.
�/�  �        �_���_�#  � +       �/@7���/�  � ,       �_�;W��_�  �        �?@&���?�  � 9       +�_�6���_�	  /� 	       W�?@���?�#  � #      
��_�k���_�  /� V      U_��@2�����  _@       ��P�4��P�  ��       ����@�����% _@ 5      ��A~�6��A�	 
�� +      ��� >���� U�        �P~�&�P����       ��� w����U�  (      T � ^T ��!���  7        �� ~  �����T  G       W� . W��Q���  q       R�� � R�����@  T      U/�� ?U/�����   �      ���` �����U    V      ���������@      �      ��� ������    �      ��� �����A    �      ��@ ������I    �      ��  �����          UP  ?�����    �          ����� �    �          =^�����    +�          K����@5    u          ����� @	    S         �����     uS         ��UU@ S0   �0         ��   x!   {i         ���   )   4��        ݽ�   "B0  rB�        4�{_  ��  +��      _����@(�9H�\      z^w�Z󕡊�����      ���{\~6���;e>���      �
�]c7�L䢜7�L䢜      �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            