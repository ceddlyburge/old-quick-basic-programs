��r�V�        ���         ���      `  ���`       ���    �   ��    �p  ��?p   �   � ;    ?�   ��1    �   ��1    ��   � !   ��   �     UP�����   ��UP�US  ��   �     ��   � !    �   ��1    ?�   ��1    �   � ;    �   ��?    �   ��        ���         ���         ���         ���   U    
��   ʪ     �   ��         �          {�          � �         s�          ��         s�          ��         #�          � �         �          ��         �          ��          �          �?�                     ���                     ���                     ���                                                                                                                       