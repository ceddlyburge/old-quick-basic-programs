��k6 d0 0 ��> FCh�߹�Ch�߹�      ������ !
E���
      _���;ޠ
�'�0���?      M�����,�%��,�%�:      k�����Ԁ B��ۯ�C      �����  �  �����      ������     �����      ?�� ��?��������      � � <`��?�������      <   p������������      �> �'�����?�����      �À�������� <  � � �� ���?��y� � � 1 ��� ������{� �  � ���������?����� a   0s� 8������������     �� G��?�������      � � =���������      > � �����������      ��?����  �����      ������,   �,��/��      |������   �����       �����X\T����]U�      7���}�� �!�hEN�e      ������ 1AE�1[      �����h"J%l+Z-+      k�����Ԁ B��ۯ�C      s���ތ  � !������      ������@    S�����      ��� �@?��O�����      _ � =���?�¿�����      �   p#�����?�����      X> �������������      �À����?���� <  � q ��� ������y� � � � �� ���?��{� �  � p������������� a   ps� 8������������     x� ���?��������      | � <����Ï�����      > � �����	������      ?�?�����  ������      S������   ����/��      ������C   C����       �?����� `���d      k������z ܜz ��      ���3��A�`�A�s�      ���^��8-��p8+-���      �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            