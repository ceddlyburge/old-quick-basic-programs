��r�ݲ0 0 )X�!$�����m���gm��� �(   �B�m?���-?�����
*D�.h F����/nߟ��.nߛ
Pj�� i؍�� ������������@G�"*e��w��v~w�}
bX0���<�o���~�N���~�@"h
1H�W����������w�ۻ���� ���C�1�����1�����q�pH�` �}��}��}��}�� �����	�"A �߿���9߷ɾ�PERB1) ��#�{u����yu��F  	� "O�.���O�.]��� �a� #���_���6+_����Q�������>˯<��>�PBb�@�ԇ��\�����T������@ CER���m��W�e�Ww��I�@@)b����o����o�Rh$ XA ��Z��6��Z��6��`��\ ����������������/s@D��čgۿ��ngۿ��L"@� Q�d��?Q��U�?Q��U2� 	� 0���v����p� ��p@�B�{y����cy����AEL� @C%2!P{����S���7�� ��� :��{�����{���?�� �`3_��Ow_��Ow�9����� ���?�����=����� $R��w���w���"�/  A�-��