�;���d0 0 �� d�2Ah� 9�Ah� 9�  d� ���$��  !
E� a
  $� _��$�ޠ"�'�0� F?  	&� M��4���,�2��,� :  6� k��4��Ԁ	��B��@ C  �� �w�0����� �@ �  �� ��_1�� ���N� ?  �� 7�1�������� �  �� �?R9_l`ؚ�0�a�� 3�  Z�@ ;s�9z��:�笀 '[  z�@ ջfig*Ds��:t  1�  w�@ ���i{� �#?s$  6  �k@ �{�Iw���1 �  < �y@ �I_��Hw  ?�`   � wi@ ����^?Ǡ�$�  � ��@ =��O����   S ���@ �����A�}��h   ����� ����}�ؔ �     ��ٽ  ���'w������   ����  �$?�0%π    ��?� <��$?��%L��    ����l� $?��L�      l� ���?��L��    ����L� >t=�?øȆ!    e?��̠ �tN.��舑A    [��Π ��B:� ?�    -+��J� ��rC;� �,	�P    ���K� ���z� ��  � ���  ��}�� A�  @ :���  ����x� �)�O   o����  g�.�{�g�ͣ`  � ,�g��  <��y�<�   �< �  �o��������� T�� /�� ���M�� �"� "  /_� z�oMf��`�^�p� �  /_@ ����|� Q�% �@ e  �@ f��N{��CϹg� �  _@ ]o�Lw����u��@ ,u  �@ ��Lo��$���v� O  �@ Y��@~� ���`� �  Y` ?t�?������A�ǀ I  }Ϡ ?���.��r���v�r� ~  }Π ]���;�P!����  �  5ހ �۔�?�@f1�� }� �  5�� �������   =� k�D;���	aܜ  �  e  ���D�A	a �A  3�  e  ��� -�8#Rp8+  {�  #  �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            