���  d0 0 < 4^���_�-� �       � �� ? ���
  @ 
      \�^���_�� �       �� 0?��p @       ��^ P�_�� �       ��=  ��?�   �        ��^��_��� �        �? ��?�	  � 	       �^���_�  �        �? ���?�	  �        �^�W��_��  �        �? ���?�  �        �^����_�   �        +�?  ���?�  �        W�^����_�   /�       ���� �����  W@       U_P~���P�   ��        ���� =�����
 w@ 
      �� ~ 7�� � ߀       ��P� +��P�� �@       �� ~ ?�� � *߀       ���� ����� UU?@        UT ~ UT � ����           � ^   ��!���@ e      UT ~ ?UT �����       ���� 4�����UU@ +      �}@^�/�}@_�
��� 1      �� � �� �� �@       ��P^���P_�  ��       ���? ���?�  W�       U_�^����_��  /�       ���? ���?�  �       UW�^����_�  �       ��? ���?�  �        W�^����_��  �        +�? 
���?�  �        �^�	W��_�  �        �? 
���?�  �        �^�U��_��  �        
�? ��?�  �        �^��_�  � 	       �� 	 ����  @        �~�_��  �       � �� @���� x @       �t^�p_�_�p �       � x� ����X @       x |^��_�_�� �       � x� 8����08 @ 8      �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            