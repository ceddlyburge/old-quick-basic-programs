�j�  d0 0 ^k��h}��ԟ������      �k���z�@D�z�@���      ����Ϡ  8�>?��9      |������p   �����      �O�����   6�����      [��UU}�  ���7�����      ��� ?� U��������      �   � ����������      �� 
� U����������      �`_�� �����������      ��+��� ����������      �_���J�����������   UT P�`~���`���`  �����  =���  ?���  ?  	�������^����_����_ W���U] W�/�� W�/�� W�/ ������ ���� ���� �� ������4����4����4�� ������V��B��V��B��V��B ����[�+��[�+��[�+��������?����?����?�������q�/�q�/�q�/�������P���7�P���7�P���7��_�����@��	��@��	��@��	������������������������������B����B����B��������W�����W�����W��������V���� ���� ���� ����/������ ����� ����� �����_�G���_�G���_�G�������U+�����+�����+���������  �T����T����T���o���  @ ���@ ���@ �������  �G���G����G���k���  �����������������T�  �����U������������  ?�  U���� ������������  �   _��� ������������  ?�   ��ª�����U������  �  ���������*������  ?�  ������U���������  �  }��������� ������  ?�  ��������� ������  �  ����� �����������  ?�  ������?�����  �  ΋����1���Z?�����  ?�  �G���� ����3�����  _�  n���������
������  ?�  �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            