���  d0 0 Hb|�=����³����      �{�_�P��� P���@      {ܿ����#@P�cSQ]      ��S�۲@Y�4M\٬4�      n��o�֑�+�J�+/      {��� �B,1� �f�1�       Z��   �`  �r�         [��   $p   /ps         |�   �   ��         ��UU@'   U�          ����� JT    �\          w���  �    �          ?���P	�    �          x�����    �      UU@ 
_�����    �      ��� �����     _      ��� ������     �      ��� _���� �     �      ����������    C      ��@ ���P��    �      ���� ������TU@   t      UU�� ^UU���!��   c       ��� v ����	�U@  )       W� | W�����          +� '  +�����  8      P � -P �����        ��
� ��
��U_�        uTz 
uT�����       ��� ����
 }  
      ��Az ��A� 
��       ���� ����� _@       ��A~ ��A�  ��       U�� 
�����  _@       
��~�����  /�        W� ����  @        +�?����?�   /�         �_@_��_�	  �        
�/�
���/�  �        �_@U��_�  �        ��

���  �        �/@��/�  �        ����  �        �/@
��/�  �       ���_��  �       �z/@@��/�` �       � ��@_��	` �        z/@�?�/� � �        � ��_�� �       �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            