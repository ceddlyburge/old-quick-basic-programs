���  d  � � � � � � � � ��������      � �     0 � �     0 � �       � �       � �        �  �        `  ` � � �    � � �    � � �      �  �   �  �   �  �        �  �        �  �        �  �    � � � �    � � �    � � �   �  � �   �      � �      � �      � �     � �    � � �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     