�j�  d0 0 ΋�˯�1���X?����\  ?�  �G��� ���3���;  �  n���������
������  ?�  G��������������  �  ����|{A�������  ?�� _G��{���迆�����  �@ ?���\=���_�����_�  ?�� ����?��������  �� _���>�_��������  ;�� ��}�/�}����}�  �� _���>���������  �� g�t�N���O����O�  �� ���_�> �_����_��  �� z�to���o����o��  �� ��:�=������  �� R|}����������  �� ��>φ?.A�χ�.��χ�  ?� }�������?���   �� ��.��?I�����M�����  � ��_L��\���   �� K��/�>��/�����/��  �� {�z�/������  �� ���>�<h_�>��o��>��  �� �E�__��_���_�  �� ?��<z>��<����<�  �� ��q�_��q�����q��  �  E�7迀��7�@���7��  �  ߢ�� _���#����  �  ���E� /������  �  ;�x�+����� �?����     ���_���������      ��O��H���� i����P      ^�R�{���������      ��@�� ���h&����x      ���_P1�7��s�      ������x>& {��6       ������_v���6_      �z��]�"���:��Ϻ�      7������"@)A�#N)C      ������h"@)Ch#N)C      7�S�y���%����-��      ��^��� �N��3?      �w����4� �u��      k�����Ԁ B��[�C      M���e��,�%��,�%�:      _���;ޠ
�'�0���?      ������ !
E���
      ��> FCh�߹�Ch�߹�      �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            