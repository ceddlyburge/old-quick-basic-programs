���  d   k  k  k  k      ~          ~  H       �     � � �� ��  �  � �  �       ?                    x  x        �  �       A� A�       c� #�       3? ?       ;��+��      ππ      ?��      ?��      ��      ;� +�       3� �       a� !�       @� @T        x        x   0 <0 <0 <0 &` 7` 7` 7` 1� 3� 3� 3� � 1� 1� 1� �  �  �  � ��������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        