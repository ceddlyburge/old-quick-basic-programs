�;��0d0 0 ��> FCh�߹�Ch�߹�      ������ !
E���
      _���;ޠ
�'�0���?      M���e��,�%��,�%�:      k�����Ԁ B��[�C      �w����4� �u��      ��^��� �N��3?      7�S�y���%����-��      �?=?�l`���p�a�����      ;s�}����G笘�g[      ջ_?g*D����:t�ȱ�      ���?�� 8�?s%���      �|����� X �X<      ��_���I� ?�i� �      ����>?	��$ɚE��      ��x���'�T�'�TS      �����C 	�k�mP��      �w�ʿ}�!5`���5`�      ?�v��w�Y�®��ٜ        ����  D"@  �        ����
"@�  .���    ������    � ��    �<���p}�\T�   ]U���    ��}� |�!   �e��    ������ 1A    1[����    ��� %   -+ �  ?>q�� >yP   �?>}p  a����z ���   �a���   ���0�    ��1�   ��x�w�!�   ��w���  ������}���`   ������  ���r�� ?�0    ����r   <dz� <"�    �� <fz  ��0���;�"  " ;�� z���楍c��^�p  � ��� ������ �4% �  e  ��� f������C&Ϲg� �  6�� ]o������7�Hu��@ lu  ?�� �ؖ���$�N�v� O  ހ Y�Ȃ�~� �ZL��`� \�  
ڀ ?h������N`A�Ǡ eI  
ހ ?������r�fv�r� ~  
� ]��*��P
���  �  
� ���*��@f�P }� X�  �� �,:���Ƥ`��� d  �� k�2����b�ܜ` O�  
�� ��貟�A,`�A  s�  
�� ��ȡ��8  Rp8+  {�  �� �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            