�;���d0 0 ���������%
���/^X      �w���K��e&o����      ������A* Pq�����      ����o�`) :�	i�q���      ������C����F�      �[��;������'���      w������@i	h�By�h      ��=;_�@R���Agz���a      �\��X �8��r��9��      ������Nf0�K��rg��      "?����Y�@FP  @��{�    �D}�}O �M��  Mڷ��    H�����F)�@q  �����(   ��h�����3:�   :����   ���W��GP�(   z?���   �E���{�x@H�   I��}��  
f�Y@���   ��S��  q5����	�   ����  ��> �`a�    i�-��  C�r6��0)Cz   �G�r<  ��8�?��Vd�x   ����~�  y�ۮ_ր��Q�    w�����  1@z��@&�fB    ��qf�v  �%�q�� E<f�8    �8�e�v  #�k��H�P    ��k��{  ���N�C�\    �]^�_�  )���;����Q�    ������  D!~���g    E��g  (J
a��c=%�    '��Zk}� � ����C[ )     �{�0��  #�Q!����r��	    �i��s�  i�6 ��eQ�
     N=m�w�� �Я�Rv�=P4    �6�~��@ !0Rf��C�h    O�/s�n� <*����2iC!	    �/>k�  i��*�� �"�    ��y���  �؎��� (    s*�ܮ� B2���n"`    sm�:� 1(�������    ������  x� ���?nA�    ����n�  .�q�ܙIȐ(+    N{���� *`�)���)0    �/�=� ��}��o%$    {e���  03D
=�I�I�P    '}y��K� J�7�5؁He�    ����@ o$���6�
    o>� �lP��F��(    i�n��� ���C��CpHX    ����S� � $ B        L��H5k �^����            ��
=�v��޳��T��  �       t������<��%�/            $�A$�" ?�̿��� `           �@�r��7�vޟu�
          d��1 w7z�o� "            #xG'�i�v)�~    �        !�$�Z     