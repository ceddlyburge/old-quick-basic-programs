�;�6d0 0 ��> FCh�߹�Ch�߹�      ������ !
E���
      _���;ޠ
�'�0���?      M���e��,�%��,�%�:      k�����Ԁ B��[�C      �w����4� �u��      ��^��� �N��3?      7�S�y���%����-��      �?=?�l`���p�a�����      ;s�}����G笘�g[      ջ_?g*D����:t�ȱ�      ���?�� 8�?s%���      �|����� X �X<      ��_���I� ?�i� �      ����>?	��$ɚE��      ��x���'�T�'�TS      �����C 	�k�mP��      �w�ʿ}�!5`���5`�      ?�v��w�Y�®��ٜ      �+��  �D   ��        ��݃��,B:��,S>      ��|����" ~��f�      �7�px ��XG����      w�7����� D���hD      �����������E     ������ h"@l+     �@y�{���X�;� �\�     ���K�� @ � >A��2�     >A೻��~ L�H�A$\�X     �$������I� ���M�      ���}�?��� ��ߎ� �     �ߎ���<  .EI��.�0     	}��Ro�h?�푣 H���     k?����x�� �:z�   z�xz�\থ�`�h^�p� �  � ����� FH% �@ e  � f��⻹�C"JϹg� �  � ]o�#����
u��p ,u  +� ��"o��$�
�v� O  *  Y��"?~� �L��`� \�  :  ?l"����`A�Ǡ eI  2  ?��3n��r�3v�r� ~  3  ]��#{�P���  �  �  ���#?�@f�P }� X�  �  �:#���9`��� d  ;  k�c����hi�ܜ` O�  k� ���b��AH��A  s�  j� ���"-�8  Rp8+  {�  "  �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            