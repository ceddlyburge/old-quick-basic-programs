�;�d0 0 ��*AFCh�#9�Ch� 9�  c  ������ �!
E� a
  � _��ջޠ�D'�0� F?  �� M������,���,� :  �� k�����Ԁ�B��@ C  �� �w�j���-� �` �  �� ��Zn�� ��N� 3?  �� 7�[&y����&��� v�  �  �?;l`�ٷp�a�� s�  �  ;s��:���G笀 g[  �  ջ\�g*D���:t� 1�  �  ��ԑ{� 5�?s%� v  �  �|�7���X �  X<  �  ��_��I� ?�i   �  �  ����>?	��$ɐ ��  �  ��.���'�T�  TS  �  �����C ��k�` ��  �  �w���}�"�`��� `�  �  ?�y��w��Y�®�ٜ  	�  �+�ۿ��B�@��  �  ������,B:�@�,S:��  �  |��j���"  �f�    `  7�����X\T����]U�      7���}�� �!�hEN�e      ������ 1AE�1[      �����h"J%l+Z-+      y�����X�JP�\�Z�      K����z�@��2�A�      ������L�HB\�Zʺ      ����x�I�"I�M�"i��      }�?���� �`� ���      ������.E .�64�      Ro��푤��������      ������ �"�"      z�_�f��`�R�^�p�[��      ����|� J�% �JE�e      f�׼���C(ÄϹg�ӌ�      ]o������Hu��{Glu      �ǿo��$�@��v�@�O      Y��߿~� �"L��`��\�      ?m�������`A�Ǿ�eI      ?�����r��v�r���~      ]�����PQ��)Q��      ���5?�@f�� }��؈      �?����� `���d      k������z ܜz ��      ���3��A�`�A�s�      ���^��8-��p8+-���      �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            