���  d0 0 � �� 8?���08 @ 8      �tz _�� �       x�� �?���� @       xt~ �_��� �       ��� @?��� h @       X�~��_��� �       8�� 	������ @       �^���_�� � 	      X�? ���?�� �       x�^���_�� �       P�? ���?�� �       p�^���_�� �       ��?  ��?�  �       p�^���_�� �       ��?  ��?�  �       P�^���_�� �       ��?  ��?�  �       p�^���_� � �       ��? @��?�'@ � '      ��^�'A�_�@ �       X� :���� @       x�^�o��_�� �       ��� 4h?���Kl @ k      ��~����A � [      ; �������a�    �      } �������   �      ~�W�������@ǀ  @      Ҹ
�/@���/�  �      �  �T�0\  9      :  ��Ŕ  )�׶  ��      ����}(  S�l S�      �����C 	�k�mP��      ��x���'�T�'�TS      ����>?	��$ɚE��      ��_���I� ?�i� �      �|����� X �X<      ���?�� 8�?s%���      ջ_?g*D����:t�ȱ�      ;s�}����G笘�g[      �?=?�l`���p�a�����      7�S�y���%����-��      ��^��� �N��3?      �w����4� �u��      k�����Ԁ B��[�C      M���e��,�%��,�%�:      _���;ޠ
�'�0���?      ������ !
E���
      ��> FCh�߹�Ch�߹�      �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            