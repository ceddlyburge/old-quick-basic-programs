��k6 d0 0 �����������            �� ���  �        �  ��~���         �� ����� �        �  �����U           �� ��~��     �   �� ���vU       �   �� ��v�      �   ��� ����vU           ��0 ��>��           ��0 ��>��U           ��� ��>���           ��� ��?��            ��� ��?���          ��� ��>�          ������>��           ��0���>���p    w     ��0���>��p    w     �����������            �����������                  ������                 ������                 ������                 0��0���1�<            ������                 ������                 ������          �����������           �����������           � 0 � >�            � 0 ��?� �< ��  � � 0 ����� �<���� ��� � 0 �ݾ� �<݁v� ݀v � 0 �˾� �<ˁ�� ˀ� � 0 ��׾� �<ׁ�� ׀� � 0 ��˾� �<ˁ�� ˀ� � 0 �ݿ��<݀�� ݀� � 0 ���� �<���� ��� � 0 ��>��<��  � � 0 �� >��< ��   � ��� ���� �< ��   � � 0 � >� �0 ��   � ��0 �� ?� �0  ��   � � � �� ?� �0  v�   v ��� � >� �0 ��   � ��0 � >� �0 ��   � � 0 � >�            �����������           �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            