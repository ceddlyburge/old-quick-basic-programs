�;�p d0 0 ��> FCh�߹�Ch�߹�      ������ !
E���
      _���;ޠ
�'�0���?      M���e��,�%��,�%�:      k�����Ԁ B��[�C      �w����4� �u��      ��^��� �N��3?      7�S�y���%����-��      �?=?�l`���p�a�����      ;s�}����G笘�g[      ջ_?g*D����:t�ȱ�      ���?�� 8�?s%���      �|����� X �X<      ��_���I� ?�i� �      ����>?	��$ɚE��      ��x���'�T�'�TS      �����C 	�k�mP��      �w�ʿ}�!5`���5`�      ?�v��w�Y�®��ٜ      �+���|�D"@���      �����,B:"�,S>.      �|���` �"  �f��       7�� ��X[�?���X     �?7���0��  3��hE@      3������� |E�     ������h"� l+@     ?ߟy�����X� y��\�      ��K���?��@�2�@     ?����� L�HG��\�Z�     �߶�����I�"A��M�"`     ��}�?�Ꮒ ���� �      ������ .E �.�64      �Ro�  푤�� �����       ������ �"�"      z�_�f��`�R�^�p�[��      ����|� J�% �JE�e      f�׼���C(ÄϹg�ӌ�      ]o������Hu��{Glu      �ǿo��$�@��v�@�O      Y��߿~� �"L��`��\�      ?m�������`A�Ǿ�eI      ?�����r��v�r���~      ]�����PQ��)Q��      ���5?�@f�� }��؈      �?����� `���d      k������z ܜz ��      ���3��A�`�A�s�      ���^��8-��p8+-���      �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            