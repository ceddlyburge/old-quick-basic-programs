�;�hd0 0 ��> FCh�߹�Ch�߹�      ������ !
E���
      _���;ޠ
�'�0���?      M���e��,�%��,�%�:      k�����Ԁ B��[�C      �w����4� �u��      ������ 
0��3?      =������?�  �?�4a 8   ������d��pd���� 1� >p1w�w���4�c��u���    c������ ��i1��� ��  ��S���~����~~��� ~ ����?�/������Y������ ���~���>����������>���_7��
O���}*���}  �|��+~��!�ԟA�%���M �  ������C�|C�c�~K��x ����[��Mէ��m���� ���;���}������ϚFۯ � ����w��'�'ɟ4     ������,B:0O,S>4O      |������"  �f��       7�����X\T����]U�      7���}�� �!�hEN�e      ������ 1AE�1[      �����h"J%l+Z-+      y�����X�JP�\�Z�      K����z�@��2�A�      ������@
Z0�ʺ      ������B?� 
C?�*0� 8   {��������?�����?� 1� 8�w�{��/�4���/�u���    1�_���w�����4����u ��  ��S���~���~�� ~ ��?�7�S����~�����~�� ~ ���?��>���������>�e�_;���O���>�����  �>^��5�_�!��O��%��� �  }������|!���~%��x �^��]���Mգ�|�m���~ ��x�������M��ϚCm� � �7��{���'���'�Ϛ    �]����ܢPX'��)Z'      ���5?�@f�� }��؈      �?����� `���d      k������z ܜz ��      ���3��A�`�A�s�      ���^��8-��p8+-���      �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            