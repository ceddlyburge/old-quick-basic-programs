�;�Pad0 0 ��,�FCh�(9�Ch� 9�  �  ����^� 	j!
E� a
  �  _���;ޠND'�0� F?  �  M������,�F�,� :  ߀ k�����ԀFB��@ C  ΀ �w�����8N �` �  ΀ ��I�� �lN� 3?  }� 7�Iy���8&��� v�  99  �?�l`��0p�a�� ��  =1  ;s����-rG笀 g[  =s  ջ1g*D�F��:t� ��  w  ��6/�� 
�?s%  �  >�  �|f{���;�X �  X<  �  ��s���H�8 ?�h  �  �x  ���>?	�=��$� �� ��  ������'T�  TS ��  ��y��C�`�k�  �� ��  �\Cz�l� E ��  � Cp  ?���!D�� � ��   ��� f?G       o����� ~  ?�9�      �����?��� <  �      �?����}� ?�}��?      �}��?����   G�~      �����x � ���~ @      ��~���  ���      ������ � ����~      ����~�q�  �| >      ���  3��@����      �3���`�`?o��  ��      p�`?�����><���9      ���=� ���8���?      ���������� ���      ������������� �� ��w�_�a��`��^�`����� ����� J�% �JDe    � f�׽���C(�DϹg���   � ]o������Hu��{Glu      �ǿo��$�@��v�@�O      Y��߿~� �"L��`��\�      ?m�������`A�Ǿ�eI      ?�����r��v�r���~      ]�����PQ��)Q��      ���5?�@f�� }��؈      �?����� `���d      k������z ܜz ��      ���3��A�`�A�s�      ���^��8-��p8+-���      �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            