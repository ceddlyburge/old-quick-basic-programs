���  d           � � � �  �  � ?� 
�  @ @ s� -@      q�        }� "@       ?�    @  @ � @  `  ` |` |`  0  0 �0 �0      A� �       c� C�       3? #?       ;����      ��K��      ?π/π      ?π/π      πKπ      ;� �       3� #�       a� A�       @�          x        x     ?  ?  ?  !` c� c� c��������� �������� � � � � � � �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         