�D�  d0 0 ^k��h}��ԟ������      ~:޳�?�šl�ؙե|��      �Z��z^0�Q��8��Q��      ���o�� �H:5�ȝ      � v��  I  �  Y  �      �                                               � *�                   UUQUU@                  �����                  _�����                  ������                  ������            *��*��������            UUUUUT������            ������������            ������������            ������������            ������������            ����������U UU       UUUUUUUUUUUU������      � �� �� �� �W�U_�U                  ������                  ������      PUP UPUP U������      ������������UUUUUU      UU��UUU��U�� *��      ������������            ������������            ������������            ������������            UUUUUT������            ��*��������                  ������                  ������                  _��_��                  ������                  UUQUU(                  ����D                  T T                     "                                   @ ~�  �     `       �
��� 8( A08� C      |�߷���t`H*�~`ʪ�      ���㿠<@�>1>l      �k���z�@D�nz�@��n      ^k��h}��ԟ������      �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            