�;���d0 0 ��> FCh�߹�Ch�߹�      ������ !
E���
      ]���΢F
3�?FQ�3      N�8�����B�   r      j�?������/�� ( #      � �����,� f&�14      �C����4�� ��      7��������	��O      � ���`}@��a�O8      ?������>��<��      �9���/��38 �@3      �   �`�Cw����'      ������e( � �(      y�s�0������� � ?      ��� ? � �� @��      ��D%��H�D��H��G      �q����@���@i � d      ��>���_�:�J�9>�      ?���?�� � �\#Z�      �+�����D"@��      ������,B:"@�,S>.��      |������"  �f��       7�����X\T����]U�      7���}�� �!�hEN�e      ������ 1AE�1[      �����h"J%l+Z-+      y�����X�JP�\�Z�      K�s�:��@(��~�G��      �/���C��?�P  �      ��_��K����J � �      t�@��3ȳ<���M���      ևhp?-���/x��      _�8�����s��<      �}��0���<�"      ���|������x"�.      �<s�:���� � �      ` > ���������      _���Z���|l��9
��      |��8ƃ��?�;� @ �      _�� ��#�?�<0�      	n��� ��	����i      >��:������  �      Q~}�߮����"��r�/      ������D0 C  v�Fk�h      �?����� `���d      k������z ܜz ��      ���3��A�`�A�s�      ���^��8-��p8+-���      �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            