�g�  d0 0 ��> FCh�߹�Ch�߹�      ������ !
E���
      _���;ޠ
�'�0���?      M���e��,�%��,�%�:      k�����Ԁ B��[�C      �w����4� �u��      ��^��� �N��3?      7�S�y���%����-��      ������h"@)Ch#N)C      7������"@)A�#N)C      �z��]�"���:��Ϻ�      ������_v���6_      ������x>& {��6       ���_P1�7��s�      ��@�� ���h&����x      ^�R�{���������      ��O��H���� i����P      ���_���������      ;�x�+����� �?����     ���E� /������  �  ߢ�� _���#����  �  E�7迀��7�@���7��  �  ��q�_��q�����q��  �  ?��<z>��<����<�  �� �E�__��_���_�  �� ���>�<h_�>��o��>��  �� {�z�/������  �� K��/�>��/�����/��  �� ��_L��\���   �� ��.��?I�����M�����  � }�������?���   �� ��>φ?.A�χ�.��χ�  ?� R|}����������  �� ��:�=������  �� z�to���o����o��  �� ���_�> �_����_��  �� g�t�N���O����O�  �� _���>���������  �� ��}�/�}����}�  �� _���>�_��������  ;�� ����?��������  �� ?���\=���_�����_�  ?�� _G��{���迆�����  �@ ����|{A�������  ?�� G��������������  �  n���������
������  ?�  �G��� ���3���;  �  ΋�˯�1���X?����\  ?�  �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            