�;�X|d0 0 �� d�2Ah� 9�Ah� 9�  d� ���$��  !
E� a
  $� _��$�ޠ"�'�0� F?  	&� M��4���,�2��,� :  6� k��4��Ԁ	��B��@ C  �� �w�0����� �@ �  �� ��_1�� ���N� ?  �� 7�1�������� �  �� �?9_l`؊�0�a�� 3�  
�@ ;s�9z���笀 '[  �@ ջFig*D���:t� 1�  �@ ���i{� #?s%� 6  k@ �|�Iw��1 �  <  y@ ��I_��I  ?�i   �  i@ ����^?	��$ɀ �  �@ ���O����  S  �@ �����C ��k�  �  �� �w٭}� � ���  �  Y�  ?�I�'w���®� �  M�  =+�$?��π�� �  _�  ��$?� BL�� S  �  Wl� ��$?� "L�  &�  � l�  �?�?HL�� 
� �? <L� ��=���Ȇ!  @ e��<̠  �N.�9��A   [8Π ���B:���    -+��J� x82B;�a�,	�P    �y�K� @��z|~ ��    �|��  ����}��    :Ǐ��  ���x��ɡO    o����  n��{�`͡`    ,�n��  ����y�~8E�    �����  �<�����<�    T��<��� � �L���"    "Ϗ^� c>Lf���^�   ��_@ ��+�|����%    e���@ fQ�N{��O�Ϲ   � _�_@ ]I�Lw����u��  ,u ��@ ��Lo��$x��p  O ��@ Y��@~�&��`  � �Y` 84�?���	��A��  I =Ϡ ?��.��q���v�p  ~ �̠ ]��;�P�����  �  �܀ �ڔ�?�@f1�� }�  �  ��� �����9���    �� k�\D;���	aܜ  �  ]e  ���D�A	a �A  3�  ]e  ��� -�8#Rp8+  {�  ~#  �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            