���  d  � � � �     �         �  �    � x �   � x � x  x  � x        � @       �  �        �  �       � �       ��      �0�       �`�@      ��Π      ���@      ?�?�      ?�?�      ?�?@      ����      �`�@      �0�       �P       �  @ @  @  @� @  `� a� a� a� 3  7` 7` 7` ` ` ` ` @ ` ` ` ( h h h � � � �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         