�;��Vd0 0 ��> FCh�߹�Ch�߹�      ������ !
E���
      _���;ޠ
�'�0���?      M���e��,�%��,�%�:      k�����Ԁ B��[�C      �w����4� �u��      ��^��� �N��3?      7�S�y���%����-��      �?=?�l`���p�a�����      ;s�}����G笘�g[      ջ_?g*D����:t�ȱ�      ���?�� 8�?s%���      �|����� X �X<      ��_���I� ?�i� �      ����>?	��$ɚE��      ��x���'�T�'�TS      �����C 	�k�mP��      �p{ʻl�% ��% �  x   ?��!D���� �8    �� �?       �?���� ~  ?�9�      �����?��� <  �      �?����}� ?�}��?      �}��?����   G�~      �����x � ���~ @      ��~���  ���      ������ � ����~      ����~�q�  �| >      ���  3��@����      �3���`�`?o��  ��      p�`?�����><���9      ���=� ���8���?      ���������� ���      ��������q����  �  � �q�w�_��%�`��^�`�  ^��� ������ J=�% �J  e   =� f��s9��C(k�Ϲg�  �   {� ]o��s����lu��z  u  �| �ā���$����v� O  �� Y����~� 顼��`� �  �� ?a�߾���% A�ǰ I  �� ?��d���r�e=v�r� ~  e� ]�����P�d��  �  �� �����@f�P }� �  �� �+)����`��� $  �@ k�)����w��ܜ` �  �� ���a��A	��A  3�  i� ���	-�84 Rp8+  {�  	  �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            