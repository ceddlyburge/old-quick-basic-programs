�;��vd0 0 �!HN�@t!     �!H@ �x���(5wh*    n�}�� �k���C    珋{�� �|���F:ԤP    �_���� ����}�� <U�    �����@ )  $��H���a    vqi���  ɚ��8� ��    O�8ͺ�  ������H �l    |��˴�  �R��}�n���A    �G����  �1��]��^��    �����  "6=2��YƆ�,    l�{���  [DM�] �[���    >�[�_�� ���_�F*J�,    s,��+�� ��h<_��_��     ����� (��w7wGP�>Ȩ    �o��� �E����x@EL    ��}�� 
e�}@����    �S��� q3�;�̀D     g��� �f ��     -��� C�r<3 0 �x      G�r<�x1�8ߙ��Voc�      3�~����y���V����      �����1@z�?@&�gp�      qf�w��e%�|a� E<b       ee�~o�#�n H�P      k��~�N�C���      ^�_����)���0���x      ������!~>|�^?�      ��~ߨJ
�Tc 0p      �Zk1� ��>C[!�      W0������Q  <]�r� �      ��s� �i�6 ��eQ�a�      m�w�����xRv�?�       W~���x!0R~ C�G�     /s�� <*����2iC/     >k���i��8� �      y��� u؎�y 8��    �wܮ�� �2C�o�    �:� �1(�oI���H�    �����` �� ��|?n �    ���n�� ��q�IȐ.�    ?ܿ��� *`�)���)��    �/�=� ����o%     5���@ 03D?�I�I��    �y��K� J�7�5؁I�*    {��� o$�;�6�    o>�  `lPקF��HX    �nn��� ��C^�CpH!H    �S��S` �߀�)	�     � /�=�  ��߀�o%      5 ���`  03D
��I�I��     � y��K�  J�7��5؁H�*     { ���  o$�;��6�      o>�   �lPק�F��HX     � nn���  ���C^��CpH!H     � S��S`  [ON���              [ON�      