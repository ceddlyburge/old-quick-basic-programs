��rȲ        ���    �p  ��p      ���    p  ���p    @  ��@   > p  ��p   |    ��    �   ��    �   ��    �4P�W�   W��0�7  ��   �    ��   �    W��0�7   �4P�W�    �   ��    �   ��    |    ��    >    ��        ��        ���        ���    �   ��         ���   ��        �         ��      �        ,    
�   ���         8          ���         p?          ���          >          ��          |          ��          x          ��          �          ��          �          ��         �          �?�                     ���                                                                                                                       