���  d0 0 ƺ��P9E'2��9E'2��      ~:޳�?�šl�ؙե|��      �Z��z^0�Q��8��Q��      �������:52�k      �޷��!I@ �%!�@ �      ��� B-  Bm@       k�=   �(ʀ  �}�        �   ��
� ���         �7�   �$U@ʬ         [�   ��?�ʦX         o��   �@�հ�h         ���    �0���(�0         z��   ��A�����P         ���*��W`1���_��         ���UUT���	          �����@���@          |_�����������          ���������ݐ�         �΃���1���1�         �����T��V U       ���UUiP��UUiR�*��      ���� �� ���_�U      �|�   (�   (� ���      u�   ��   �����      {
�P U��P U�� ���      O���������වUUU      ����U�U *��      }����������M�         ������������          o����������ك          ]������A�����          /��UUTу���у@         N�પ��"����         �4�    �C���a�@         ?{�   ��1�����0         i��   ��P_�ꟻP         o��   � *�՘0         ޯ�   )QU(-S�         ���   @��@;��         ?��   �B`T ��r         ]7�  ���   ���         �ڠ  ��%�  �ӭ�        [���  � 6D       �J��߶�8($I6�8�$k      |�߷���t`H*�~`ʪ�      ���㿠<@�>1>l      �k���z�@D�nz�@��n      ^k��h}��ԟ������      �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            