�;�@�d0 0 ��> F2Ci�߹�Ch�߹�      ������ !
E���
      _���;ܠѪ�/����?      O��e��-����-н�:      ;����ԇ�B��[��C      �s����5�$�u��      ������   �3?��   ?���Y6� ��� �����   �{�2�, ����  ���?��   z{�}�懇��G�  �g[��   ���?�d  ���   �����   �������H?   j����  ������	   X"   X>���  ��?�����(q?   zq����  ������   ��   E����   9��h���?�T�� �T�?��   �����@ 	P�` P����   �����u  '4 �  '4 ���� =}~��g� <�®�� �   � y-�����d |��    ��������?<f'��<w     ���|������#���g�    ?���wÏ����<~< ��     ���7������ @��h     ����������ǀyE     �����������   	l�     ����5������� >��     ����K������������    ���;;������@�|�@    ����^����M�`  M�`    ���}�.���� �t� ���      ������.   6.�  7� ?��  �o��?��� �� ��  e����ߚ  >�   ����� �������^�   ����� ����ڀ~�s%    e?���� ~?���0�� ~ π    �?���� o������   u�   u���� ��������     O���� ���o� ��    ����� ������ � � �    ����� _���ꋿ� �v�   ~?���� �������  ��?���  ����?�@ Z�|  ^؞���  _�����  `R��	d^ �   go����ܐ~0-ܜ~0��      ���7M��`�M��s�      ���^� -��h ;-���      ꋀ�� �v �   ~ ����  �������   ���?���   ?���?��� Z� �  ^؞ ����   _�����  `R���	d^� �    go�����ܐ~0- ܜ~0��        ��7����`� M��s�        ��^ퟀ�-��h  ;-���        ������� �2� � �2�            