���  d0 0 n���������
������  ?�  �G���� ����3�����  _�  ΋����1���Z?�����  ?�  ������?�����  �  ����� �����������  ?�  ��������� ������  �  }��������� ������  ?�  ������U���������  �  ���������*������  ?�   ��ª�����U������  �   _��� ������������  ?�  U���� ������������  �  �����U������������  ?�  �����������������T�  �G���G����G���k���  @ ���@ ���@ �������  �T����T����T���o���  +�����+�����+���������  _�G���_�G���_�G�������U����� ����� ����� ��������� ���� ���� ����/��W�����W�����W��������V���B����B����B����������������������������@��	��@��	��@��	�������P���7�P���7�P���7��_����q�/�q�/�q�/��������?����?����?�������[�+��[�+��[�+���������V��B��V��B��V��B ������4����4����4�� ������ ���� ���� �� ����U] W�/�� W�/�� W�/ ���Ъ���^����_����_ W�����  =���  ?���  ?  	���P�`~���`���`  ����_���J�����������   UT ��+��� ����������      �`_�� �����������      �� 
� U����������      �   � ����������      ��� ?� U��������      [��UU}�  ���7�����      �O�����   6�����      |������p   �����      ����Ϡ  8�>?��9      �k���z�@D�z�@���      ^k��h}��ԟ������      �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            