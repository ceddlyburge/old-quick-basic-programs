�;���d0 0 ���E�K/ �<����      ��_��)��0$�}��q$      ��[FΎ��3q����w�      ������Fm#K���/c[      v����\�Y��^���      ����{�1�(�";�����      �����+T�0�?�����      ��v���@*�`bu������      ݯ�����P���  z  �� _����Ix\���  � ��� {v=4[��������  � ��� ��M�m�D[��WWP  
w _�� ���+2&*D���  � +�� �4h7w���Z 7�  � �p ��s#ߤP�=� ��  a ;�� �Ű�&�%x@9e�  = }��< u
d�������  � E�� ��q7��-���   � ��� ψ�#�8bO~�   �$ ��r4���0(B��  � gr<� ��8��& �Vg2�#�  � c~�� ���ۃ~���<�߀  � y��� �@z�%��g���  � f�w ���p3�E<f!-�  ' e�v0 ��kZ�x�P�h}�  n C�{� ��ӽ@BC��BI   � __�� �)��� ���@h�  r )�� ޡ~�%�g0T-�   T ag0 ��
a�{2�c=n�s�  � Zk}� � ����Q�[ 6�߀  � 0��� �cQ!��0�r��P��  ~ ?s�� �u6 ���Q�Q��  u w�� �����=�!Y�  � ��� ?�Rf���C�h	/�@  	� �n� Kڬ��ߵ�C!08��  } ﳰ }��*'����Q��  � �� �z����� ((��  9�  �� �����=.�)�~}q���      ��{�����PJ���SJ�      �����@h��������      Sߟ_��� p�B�����z      _M5n�}���j�������      ���߀�� �J�׻{      ۻ�w��e������_      �{����-�Cm߯*[U      ��ǝ���xb���|��a      ~�����r����{���      ߟ;�kl(���շ������      � $ B        L��H5k �^����            ��
=�v��޳��T��  �       t������<��%�/            $�A$�" ?�̿��� `           �@�r��7�vޟu�
          d��1 w7z�o� "            #xG'�i�v)�~    �        !�$�Z     