�j�  d0 0 ƺ��P9E'2��9E'2��      ~:޳�?�šl�ؙե|��      �Z��z^0�Q��8��Q��      ���o�� �H:5�ȝ      ����w�!Im�%!�}�      ���F^� BX���BX��      ��+ݺ� �#E ���3Gh      �;��U�������X      ���{�@�������       W���]��)(�����/�       ������D#X���];Y        ��{��� 0�d���0�d      ��+������$ ����D      �P�����������      ��������@Q������      ��Po��������������      ����w����c�������      ���������QL�����L      UT��ԺUT��+EUT���媫@     �C�i  ���  ������      /���  /�?�  /������   ����������������   ����y������������   ���t�����Ea����i����  ��@����@�����@������   U�y�U��rU��r����   ?��>� ?���A ?���E���@   �]� �_�r �_�s����  U�./�U�/�U�/�R����  ��z���z���z� ?��  ��������P����Z _��  ��~�^��~����~��� 7��  ��?���?�Q��?�u ��  ��_�l��_����_��� ��  E|?�}��?����?�� ��   �������Q����s ��  `\Ϗ�����D����U ��  �.�����d����� ��  ��Ϗ����������  �  �G�� �G��D��G���  ��  �ώ߀����"�����7  �  �Ǉ\�Ǉ���Ǉ��  ?�  _ÃϏ��?���c7����c  �  ���� ?��I7���k  �  ��Ϗ��?���������  ?�  ������@����l  �  ��Ϗ�p����n����n  ?�  ^�}����������  �  �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            