�;��[d0 0 ��> FCh�߹�Ch�߹�      ������ !
E���
      _���;ޠ
�'�0���?      M���e��,�%��,�%�:      k�����Ԁ B��[�C      �w����4� �u��      ��^��� �N��3?      7�S�y���%����-��      �?=?�l`���p�a�����      ;s�}����G笘�g[      ջ_?g*D����:t�ȱ�      ���?�� 8�?s%���      �|����� X �X<      ��_���I� ?�i� �      ����>?	��$ɚE��      ��x���'�T�'�TS      �����C 	�k�mP��      �p{ʻl�% ��% �  x   ?��!D���� �8    �� �?       �?���� ~  ?�9�      �����?��� <  �      �?����}� ?�}��?      �}��?����   G�~      �����x � ���~ @      ��~���  ���      ������ � ����~      ����~�q�  �| >      ���  3��@����      �3���`�`?o��  ��      p�`?�����><���9      ���=� ���8���?      ���������� ���      ��������p����   �t��w�8�a��c���^�` ����� ����  ���% � e ��� f��ѫ��@6`DϹ`  � ��� ]n"H�����Hu��  lu  3�  �0`o��$8���v  �O  8�  Y��$�~� ��L��`� \�  �  ?L$�����n`A�ǀ eI  n  ?��fn��r�.v�r� ~  n  ]��&{�P
��  �  .  ���"?�@f�� }� X�  �� �6n�������� d  � k��{���hÍܜ` O�  � �����A���A  s�  �� ��ڨ-�8(�Rp8+  {�  �  �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            