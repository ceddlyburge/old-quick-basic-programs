��k6 d0 0 ��?��Ch�FCh�F      ����W�  (BU��B   � _�����   W�2�єW 0 � Mk�k_����d�ѝ�� � � k�w]{�Ԁ
� Z��ۧ�� r�� �7���
�T@ ��~��R�"� �����  � 
���/S@2� 5�ӭ���
 @Q���~�iU��`��,��l`� Fa�������;_�����   ����� �p��߿����    >}���7u�C� ����     w������>�����;���     ���4�{� ������ � ������ ����������    /����~ � \���� ' 8�����;ـn� ���ƾ�A  H����h|�� �煯=  8 
�����8Gq�/���� �ӿ؝����X��3����DD""%����u� H ��\���(@+BP/{�{��)�L |�����  �o�X(�	F }w���� ���ڟ^�H�F 7������  @ �iDKJ- H @ ���_���(!M�h+   @ �����Th"A�l+aX�      |�>�.}�h�т�h�у      ����� 
�U���     ������` 
@ z2��e 0  ` �k����r�ds��g}� � d k�v�^픀) ���i� r� � �7�n�
�����R��@{�~w|�� ����寿�S@������i�
 @����U��^�-��[��@����C���n8�_����$  H /��_�� �p��_�����  � �}����u�� o������    ���o��>/||p�;��v�   	��������^������ b ������ ����?����� � ������~ � \<��� '� N�����Nـ� x��񯭁 	 �����|�,����ak�G � O����v�8�po�~���� �ӿ�'��!V03��gw�DD�����?��� R ��]-�(@*ЀU/{���})�S ���y�? �@o���(�Q��� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            