�;�0�d0 0 �!H[�@t! f    f�!HP �x�ϰ(5w`O    O�}�� �k����!    /��{�� �|��F:Ԥ#�    �_���� ����O�� <Q2�    �����p )  $��H���R�    �i����  ɚ ޻8� �!�    �8ͺ�� ���w�H �4�    ��˴�0 �R����n���    <����� �1����xo    #���� "6=4[�YƆ��    {���� [DM�g� �[��     
[�_�� ����F*D�     ���+�� ��h7v���Z	    ����p (��s*7GP�=��    �o��� �E��*�x@5    �}��0 
d��@��Ԁ    �S��� q7�w���    ���� �)� �b!    1-��  C�r4��0(<    �G�r<� 1�8����Vg%'    '3�~�� �y�ۘ�V���/    ������ 1@z�@&�gH    Hqf�w  e%�p?� E<f K     [ee�v  #�ky�H�P�    ]k��{� ���N�C���    �^�_�� �)��_}0��� �    "�����  �!~d��gD    d��g  �J
a��Tc=     -�Zk}   ����C[ (P    *�W0��  ��Q'�g]�r�b�   ���s�  i�6~�eQ��:   �:m�w�  ���Rv�%m   }W~��  !0R��C�WF�   ޚ/s�@  <*��sw2iC	��   ��>k�  �����uP t��@  v��9��   ;@�ۥ�ļ1$Z ĸ%[A �   N��������      ��w���""�Ws&2�RWw      ������wX3�wx�ڶ�      ��_�<qX���q[��>�      ^���=z�!t�Ǐ�+|��      ?�����р .�H݁b�x      ���L�A ,����      v���θ�;�77g�;�??g      筽���RBb:�o�b      ��:Z���ŭnL�����      ���7�1 �؇�@����      =z��!t�Ǐ �+|��        ?������р .�H ݁b�x        ��L�A��,��� �        v���θ��;�77g �;�??g        g�������RBb :�o�b        {�:Z�����ŭnL ����� �      ��7�1���؇� ����� �      ������                         