�;��d0 0 ������      ��<�      ���S�� ��X<��;      ������ �\s�T�\�      ����g{P X��P�ڐ��      �ϴ���b0Ki0b0�i0�      o������5���5|�      o���Ͼ�!5 �A�+}��      _������z h�z	��K      }��﷗�-�hǨ?��h      o������@    ��         &&?w9zYڄ�ƀ� �ƀ@�  \�M�3[��D@ h� P_�w���� F*@*P  ( ��+�W��h7�9��Z   � ���~u?(��s#GP�=�X      o���Z�E��%a�x@8      �}��=c
d��@���      S����q7����*      �����# �bH      -��'MC�r4��0(*      G�r<��1�8���Vg0�      3�~����y�ۀ�V���>A      ������1@z�@&�g       qf�w�e%�p2F E<f(      ee�v3n#�kY]H�P��      k��{����0N�C��      ^�_��5�)���0���$      ������!~��g3	      ��g3٨J
a��Tc=m�      �Zk}�� ���LC[ 42      W0���~��Q!��]�r��\      ��s���i�6 �eQ��      m�w�����Rv�=�      W~����!0Rf��C�h'      /s�n��<*����2iC!1      >kﳵ�i��*� ��h      y����u؎΂K (M�      wܮ����2�n
�      �:���1(��4I���Y[      ������� �/�?no      ��n�?��q��IȐj�      ������*`�)���){      /�=����d7�o%!      ���g703D
I�I�D      y��K�^J�7�5؁H�K      ����o$�8�6�b      o>�>�`lP�F��N+      nn���/��CBLCpH8�      S��Sz�����){        /�=�����d7 �o%!        ���g7 03D
�I�I�D        y��K�^�J�7� 5؁H�K        ���� o$�8��6�b        o>�>��lP��F��N+        nn���/����CBL CpH8�        S��Sz� X�t�ǀ              X�t�ǀ    