���  d0 0 ��> FCh�߹�Ch�߹�      ������ !
E���
      _���;ޠ
�'�0���?      M���e��,�5��,�5�:      k���vԀH���[RH�      �wϽހ�4B! �uf+       ��Z�@  �   N��@       7��   �$   ��         �>�   `�@   a�`         ;w@   䈀����         խ    *R )UU:W          ��      ���s          �h    �
����          �    �%���X          �P ���W���%�          � UU� ������          �� +��A_���i           �� ��� ����           ?�������          � ���
����          � ��U*���U.   �      z ���������   UU      n �U ���U �  ��      > � ��� �  �      � /�  ��    +��      � _� 
h/�� 
h  W��      x ?PU�_�PU�  ���      P ^�*��/��*�� �Q      � ?AW�P_�AW�P  ��       � ^���@?����X }P       p ������� ��       � ~��� ����  }        P �������� �        �~�P��� �        p �� ������ �        ���  ���  �        `�� ������ �        P�P ����� �        p�� ������ �        P�/@ ��/�P� �        �� ��� � �        0�/@ ��/��� �        P�_� ���_�@� �        ��?@@�?��p �        p�^���_�� �       `�? ��?�� �       ��^� ��_�  �       ��? 0�?�0 �       �� �r��v��r���~�       ]���� �PQ‪�)Q���       ��5?���f��  ���؈ �      �?��� �� `����d�       k���� ��z �ܜz �ƀ       {��3�� �A�`�A�s��       G��^����-��p 8+-���        ^?�e�!�a�w !�a�w            